// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 18 2025 23:48:51

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_g,
    T01,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_g;
    output T01;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__50616;
    wire N__50615;
    wire N__50614;
    wire N__50605;
    wire N__50604;
    wire N__50603;
    wire N__50596;
    wire N__50595;
    wire N__50594;
    wire N__50587;
    wire N__50586;
    wire N__50585;
    wire N__50578;
    wire N__50577;
    wire N__50576;
    wire N__50569;
    wire N__50568;
    wire N__50567;
    wire N__50560;
    wire N__50559;
    wire N__50558;
    wire N__50551;
    wire N__50550;
    wire N__50549;
    wire N__50542;
    wire N__50541;
    wire N__50540;
    wire N__50533;
    wire N__50532;
    wire N__50531;
    wire N__50524;
    wire N__50523;
    wire N__50522;
    wire N__50515;
    wire N__50514;
    wire N__50513;
    wire N__50506;
    wire N__50505;
    wire N__50504;
    wire N__50497;
    wire N__50496;
    wire N__50495;
    wire N__50488;
    wire N__50487;
    wire N__50486;
    wire N__50479;
    wire N__50478;
    wire N__50477;
    wire N__50470;
    wire N__50469;
    wire N__50468;
    wire N__50451;
    wire N__50448;
    wire N__50447;
    wire N__50444;
    wire N__50441;
    wire N__50436;
    wire N__50433;
    wire N__50430;
    wire N__50427;
    wire N__50424;
    wire N__50421;
    wire N__50420;
    wire N__50417;
    wire N__50416;
    wire N__50413;
    wire N__50410;
    wire N__50407;
    wire N__50400;
    wire N__50399;
    wire N__50396;
    wire N__50395;
    wire N__50394;
    wire N__50393;
    wire N__50392;
    wire N__50391;
    wire N__50390;
    wire N__50387;
    wire N__50386;
    wire N__50385;
    wire N__50384;
    wire N__50383;
    wire N__50376;
    wire N__50371;
    wire N__50368;
    wire N__50363;
    wire N__50360;
    wire N__50359;
    wire N__50356;
    wire N__50353;
    wire N__50350;
    wire N__50349;
    wire N__50348;
    wire N__50345;
    wire N__50342;
    wire N__50337;
    wire N__50334;
    wire N__50331;
    wire N__50326;
    wire N__50319;
    wire N__50316;
    wire N__50309;
    wire N__50306;
    wire N__50295;
    wire N__50292;
    wire N__50289;
    wire N__50286;
    wire N__50285;
    wire N__50284;
    wire N__50281;
    wire N__50280;
    wire N__50279;
    wire N__50278;
    wire N__50277;
    wire N__50276;
    wire N__50273;
    wire N__50270;
    wire N__50267;
    wire N__50264;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50260;
    wire N__50259;
    wire N__50252;
    wire N__50251;
    wire N__50250;
    wire N__50249;
    wire N__50248;
    wire N__50247;
    wire N__50246;
    wire N__50245;
    wire N__50244;
    wire N__50243;
    wire N__50242;
    wire N__50241;
    wire N__50240;
    wire N__50239;
    wire N__50238;
    wire N__50237;
    wire N__50234;
    wire N__50231;
    wire N__50226;
    wire N__50223;
    wire N__50214;
    wire N__50211;
    wire N__50208;
    wire N__50201;
    wire N__50192;
    wire N__50183;
    wire N__50174;
    wire N__50171;
    wire N__50170;
    wire N__50167;
    wire N__50164;
    wire N__50163;
    wire N__50162;
    wire N__50161;
    wire N__50160;
    wire N__50159;
    wire N__50158;
    wire N__50157;
    wire N__50156;
    wire N__50153;
    wire N__50150;
    wire N__50137;
    wire N__50134;
    wire N__50131;
    wire N__50126;
    wire N__50117;
    wire N__50108;
    wire N__50101;
    wire N__50098;
    wire N__50087;
    wire N__50082;
    wire N__50081;
    wire N__50078;
    wire N__50075;
    wire N__50074;
    wire N__50071;
    wire N__50068;
    wire N__50065;
    wire N__50058;
    wire N__50055;
    wire N__50054;
    wire N__50051;
    wire N__50048;
    wire N__50045;
    wire N__50042;
    wire N__50037;
    wire N__50036;
    wire N__50033;
    wire N__50030;
    wire N__50029;
    wire N__50026;
    wire N__50023;
    wire N__50020;
    wire N__50013;
    wire N__50010;
    wire N__50009;
    wire N__50008;
    wire N__50005;
    wire N__50000;
    wire N__49997;
    wire N__49994;
    wire N__49989;
    wire N__49988;
    wire N__49987;
    wire N__49986;
    wire N__49985;
    wire N__49974;
    wire N__49971;
    wire N__49968;
    wire N__49967;
    wire N__49964;
    wire N__49963;
    wire N__49962;
    wire N__49961;
    wire N__49958;
    wire N__49955;
    wire N__49952;
    wire N__49951;
    wire N__49948;
    wire N__49943;
    wire N__49940;
    wire N__49937;
    wire N__49934;
    wire N__49931;
    wire N__49928;
    wire N__49925;
    wire N__49922;
    wire N__49919;
    wire N__49912;
    wire N__49905;
    wire N__49904;
    wire N__49901;
    wire N__49900;
    wire N__49897;
    wire N__49894;
    wire N__49893;
    wire N__49890;
    wire N__49889;
    wire N__49888;
    wire N__49887;
    wire N__49886;
    wire N__49883;
    wire N__49880;
    wire N__49877;
    wire N__49876;
    wire N__49875;
    wire N__49874;
    wire N__49871;
    wire N__49866;
    wire N__49865;
    wire N__49864;
    wire N__49863;
    wire N__49862;
    wire N__49861;
    wire N__49860;
    wire N__49857;
    wire N__49854;
    wire N__49849;
    wire N__49846;
    wire N__49845;
    wire N__49842;
    wire N__49841;
    wire N__49840;
    wire N__49839;
    wire N__49836;
    wire N__49833;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49821;
    wire N__49820;
    wire N__49819;
    wire N__49818;
    wire N__49817;
    wire N__49816;
    wire N__49815;
    wire N__49814;
    wire N__49813;
    wire N__49806;
    wire N__49801;
    wire N__49798;
    wire N__49795;
    wire N__49792;
    wire N__49783;
    wire N__49778;
    wire N__49775;
    wire N__49772;
    wire N__49761;
    wire N__49758;
    wire N__49755;
    wire N__49746;
    wire N__49743;
    wire N__49716;
    wire N__49715;
    wire N__49712;
    wire N__49711;
    wire N__49710;
    wire N__49709;
    wire N__49706;
    wire N__49705;
    wire N__49702;
    wire N__49701;
    wire N__49700;
    wire N__49697;
    wire N__49696;
    wire N__49693;
    wire N__49692;
    wire N__49691;
    wire N__49690;
    wire N__49687;
    wire N__49686;
    wire N__49685;
    wire N__49684;
    wire N__49683;
    wire N__49682;
    wire N__49681;
    wire N__49680;
    wire N__49679;
    wire N__49678;
    wire N__49675;
    wire N__49672;
    wire N__49669;
    wire N__49666;
    wire N__49663;
    wire N__49650;
    wire N__49645;
    wire N__49634;
    wire N__49627;
    wire N__49608;
    wire N__49607;
    wire N__49606;
    wire N__49603;
    wire N__49600;
    wire N__49599;
    wire N__49598;
    wire N__49597;
    wire N__49596;
    wire N__49589;
    wire N__49586;
    wire N__49585;
    wire N__49584;
    wire N__49583;
    wire N__49582;
    wire N__49581;
    wire N__49580;
    wire N__49579;
    wire N__49578;
    wire N__49577;
    wire N__49576;
    wire N__49575;
    wire N__49574;
    wire N__49571;
    wire N__49568;
    wire N__49567;
    wire N__49566;
    wire N__49565;
    wire N__49564;
    wire N__49561;
    wire N__49558;
    wire N__49545;
    wire N__49542;
    wire N__49539;
    wire N__49538;
    wire N__49537;
    wire N__49534;
    wire N__49527;
    wire N__49524;
    wire N__49517;
    wire N__49510;
    wire N__49507;
    wire N__49502;
    wire N__49499;
    wire N__49498;
    wire N__49491;
    wire N__49486;
    wire N__49483;
    wire N__49480;
    wire N__49475;
    wire N__49470;
    wire N__49469;
    wire N__49468;
    wire N__49467;
    wire N__49466;
    wire N__49465;
    wire N__49464;
    wire N__49461;
    wire N__49460;
    wire N__49459;
    wire N__49458;
    wire N__49455;
    wire N__49452;
    wire N__49451;
    wire N__49446;
    wire N__49441;
    wire N__49432;
    wire N__49427;
    wire N__49424;
    wire N__49421;
    wire N__49416;
    wire N__49411;
    wire N__49408;
    wire N__49401;
    wire N__49398;
    wire N__49383;
    wire N__49382;
    wire N__49381;
    wire N__49378;
    wire N__49375;
    wire N__49374;
    wire N__49373;
    wire N__49372;
    wire N__49369;
    wire N__49368;
    wire N__49367;
    wire N__49366;
    wire N__49365;
    wire N__49364;
    wire N__49361;
    wire N__49358;
    wire N__49351;
    wire N__49348;
    wire N__49343;
    wire N__49336;
    wire N__49331;
    wire N__49326;
    wire N__49317;
    wire N__49316;
    wire N__49315;
    wire N__49312;
    wire N__49309;
    wire N__49306;
    wire N__49299;
    wire N__49298;
    wire N__49295;
    wire N__49292;
    wire N__49289;
    wire N__49284;
    wire N__49281;
    wire N__49280;
    wire N__49277;
    wire N__49274;
    wire N__49271;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49257;
    wire N__49254;
    wire N__49251;
    wire N__49250;
    wire N__49249;
    wire N__49248;
    wire N__49247;
    wire N__49246;
    wire N__49245;
    wire N__49244;
    wire N__49243;
    wire N__49242;
    wire N__49241;
    wire N__49240;
    wire N__49239;
    wire N__49238;
    wire N__49237;
    wire N__49236;
    wire N__49235;
    wire N__49234;
    wire N__49233;
    wire N__49232;
    wire N__49231;
    wire N__49230;
    wire N__49229;
    wire N__49228;
    wire N__49227;
    wire N__49226;
    wire N__49225;
    wire N__49224;
    wire N__49223;
    wire N__49222;
    wire N__49221;
    wire N__49220;
    wire N__49219;
    wire N__49218;
    wire N__49217;
    wire N__49216;
    wire N__49215;
    wire N__49214;
    wire N__49213;
    wire N__49212;
    wire N__49211;
    wire N__49210;
    wire N__49209;
    wire N__49208;
    wire N__49207;
    wire N__49206;
    wire N__49205;
    wire N__49204;
    wire N__49203;
    wire N__49202;
    wire N__49201;
    wire N__49200;
    wire N__49199;
    wire N__49198;
    wire N__49197;
    wire N__49196;
    wire N__49195;
    wire N__49194;
    wire N__49193;
    wire N__49192;
    wire N__49191;
    wire N__49190;
    wire N__49189;
    wire N__49188;
    wire N__49187;
    wire N__49186;
    wire N__49185;
    wire N__49184;
    wire N__49183;
    wire N__49182;
    wire N__49181;
    wire N__49180;
    wire N__49179;
    wire N__49178;
    wire N__49177;
    wire N__49176;
    wire N__49175;
    wire N__49174;
    wire N__49173;
    wire N__49172;
    wire N__49171;
    wire N__49170;
    wire N__49169;
    wire N__49168;
    wire N__49167;
    wire N__49166;
    wire N__49165;
    wire N__49164;
    wire N__49163;
    wire N__49162;
    wire N__49161;
    wire N__49160;
    wire N__49159;
    wire N__49158;
    wire N__49157;
    wire N__49156;
    wire N__49155;
    wire N__49154;
    wire N__49153;
    wire N__49152;
    wire N__49151;
    wire N__49150;
    wire N__49149;
    wire N__49148;
    wire N__49147;
    wire N__49146;
    wire N__49145;
    wire N__49144;
    wire N__49143;
    wire N__49142;
    wire N__49141;
    wire N__49140;
    wire N__49139;
    wire N__49138;
    wire N__49137;
    wire N__49136;
    wire N__49135;
    wire N__49134;
    wire N__49133;
    wire N__49132;
    wire N__49131;
    wire N__49130;
    wire N__49129;
    wire N__49128;
    wire N__49127;
    wire N__49126;
    wire N__49125;
    wire N__49124;
    wire N__49123;
    wire N__49122;
    wire N__49121;
    wire N__49120;
    wire N__49119;
    wire N__49118;
    wire N__49117;
    wire N__49116;
    wire N__49115;
    wire N__49114;
    wire N__49113;
    wire N__49112;
    wire N__49111;
    wire N__49110;
    wire N__48825;
    wire N__48822;
    wire N__48821;
    wire N__48820;
    wire N__48819;
    wire N__48816;
    wire N__48815;
    wire N__48814;
    wire N__48813;
    wire N__48812;
    wire N__48811;
    wire N__48808;
    wire N__48807;
    wire N__48806;
    wire N__48805;
    wire N__48804;
    wire N__48803;
    wire N__48802;
    wire N__48801;
    wire N__48798;
    wire N__48795;
    wire N__48792;
    wire N__48783;
    wire N__48780;
    wire N__48777;
    wire N__48770;
    wire N__48767;
    wire N__48764;
    wire N__48763;
    wire N__48762;
    wire N__48761;
    wire N__48760;
    wire N__48759;
    wire N__48758;
    wire N__48757;
    wire N__48756;
    wire N__48755;
    wire N__48754;
    wire N__48753;
    wire N__48752;
    wire N__48751;
    wire N__48750;
    wire N__48749;
    wire N__48748;
    wire N__48747;
    wire N__48746;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48727;
    wire N__48722;
    wire N__48717;
    wire N__48714;
    wire N__48705;
    wire N__48696;
    wire N__48689;
    wire N__48680;
    wire N__48671;
    wire N__48670;
    wire N__48669;
    wire N__48668;
    wire N__48667;
    wire N__48666;
    wire N__48663;
    wire N__48660;
    wire N__48655;
    wire N__48652;
    wire N__48645;
    wire N__48638;
    wire N__48631;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48611;
    wire N__48602;
    wire N__48591;
    wire N__48590;
    wire N__48589;
    wire N__48588;
    wire N__48587;
    wire N__48586;
    wire N__48585;
    wire N__48584;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48546;
    wire N__48545;
    wire N__48544;
    wire N__48543;
    wire N__48542;
    wire N__48541;
    wire N__48540;
    wire N__48539;
    wire N__48538;
    wire N__48537;
    wire N__48536;
    wire N__48535;
    wire N__48534;
    wire N__48533;
    wire N__48532;
    wire N__48531;
    wire N__48530;
    wire N__48529;
    wire N__48528;
    wire N__48527;
    wire N__48526;
    wire N__48525;
    wire N__48524;
    wire N__48523;
    wire N__48522;
    wire N__48521;
    wire N__48520;
    wire N__48519;
    wire N__48518;
    wire N__48517;
    wire N__48516;
    wire N__48515;
    wire N__48514;
    wire N__48513;
    wire N__48512;
    wire N__48511;
    wire N__48510;
    wire N__48509;
    wire N__48508;
    wire N__48507;
    wire N__48506;
    wire N__48505;
    wire N__48504;
    wire N__48501;
    wire N__48500;
    wire N__48499;
    wire N__48498;
    wire N__48497;
    wire N__48496;
    wire N__48495;
    wire N__48494;
    wire N__48493;
    wire N__48492;
    wire N__48489;
    wire N__48488;
    wire N__48487;
    wire N__48486;
    wire N__48485;
    wire N__48484;
    wire N__48483;
    wire N__48482;
    wire N__48481;
    wire N__48480;
    wire N__48479;
    wire N__48478;
    wire N__48477;
    wire N__48476;
    wire N__48475;
    wire N__48474;
    wire N__48473;
    wire N__48472;
    wire N__48471;
    wire N__48470;
    wire N__48469;
    wire N__48468;
    wire N__48467;
    wire N__48466;
    wire N__48465;
    wire N__48464;
    wire N__48463;
    wire N__48462;
    wire N__48461;
    wire N__48460;
    wire N__48459;
    wire N__48458;
    wire N__48457;
    wire N__48456;
    wire N__48455;
    wire N__48454;
    wire N__48453;
    wire N__48450;
    wire N__48449;
    wire N__48448;
    wire N__48447;
    wire N__48446;
    wire N__48445;
    wire N__48444;
    wire N__48443;
    wire N__48442;
    wire N__48441;
    wire N__48438;
    wire N__48437;
    wire N__48436;
    wire N__48435;
    wire N__48434;
    wire N__48433;
    wire N__48432;
    wire N__48431;
    wire N__48430;
    wire N__48429;
    wire N__48428;
    wire N__48427;
    wire N__48426;
    wire N__48423;
    wire N__48422;
    wire N__48421;
    wire N__48420;
    wire N__48419;
    wire N__48418;
    wire N__48417;
    wire N__48416;
    wire N__48415;
    wire N__48414;
    wire N__48413;
    wire N__48412;
    wire N__48409;
    wire N__48408;
    wire N__48407;
    wire N__48406;
    wire N__48405;
    wire N__48404;
    wire N__48403;
    wire N__48402;
    wire N__48401;
    wire N__48400;
    wire N__48399;
    wire N__48398;
    wire N__48397;
    wire N__48396;
    wire N__48395;
    wire N__48394;
    wire N__48393;
    wire N__48392;
    wire N__48391;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48089;
    wire N__48088;
    wire N__48087;
    wire N__48086;
    wire N__48085;
    wire N__48084;
    wire N__48083;
    wire N__48082;
    wire N__48081;
    wire N__48080;
    wire N__48079;
    wire N__48078;
    wire N__48077;
    wire N__48076;
    wire N__48075;
    wire N__48074;
    wire N__48073;
    wire N__48072;
    wire N__48071;
    wire N__48070;
    wire N__48069;
    wire N__48068;
    wire N__48067;
    wire N__48066;
    wire N__48065;
    wire N__48064;
    wire N__48063;
    wire N__48062;
    wire N__48061;
    wire N__48052;
    wire N__48043;
    wire N__48038;
    wire N__48029;
    wire N__48020;
    wire N__48011;
    wire N__48002;
    wire N__47993;
    wire N__47990;
    wire N__47987;
    wire N__47974;
    wire N__47971;
    wire N__47966;
    wire N__47961;
    wire N__47958;
    wire N__47957;
    wire N__47954;
    wire N__47951;
    wire N__47946;
    wire N__47945;
    wire N__47944;
    wire N__47941;
    wire N__47938;
    wire N__47935;
    wire N__47934;
    wire N__47929;
    wire N__47926;
    wire N__47923;
    wire N__47920;
    wire N__47915;
    wire N__47910;
    wire N__47907;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47897;
    wire N__47894;
    wire N__47891;
    wire N__47886;
    wire N__47885;
    wire N__47882;
    wire N__47881;
    wire N__47878;
    wire N__47875;
    wire N__47872;
    wire N__47871;
    wire N__47868;
    wire N__47863;
    wire N__47860;
    wire N__47857;
    wire N__47854;
    wire N__47847;
    wire N__47846;
    wire N__47843;
    wire N__47842;
    wire N__47841;
    wire N__47838;
    wire N__47835;
    wire N__47832;
    wire N__47829;
    wire N__47828;
    wire N__47827;
    wire N__47826;
    wire N__47823;
    wire N__47822;
    wire N__47819;
    wire N__47814;
    wire N__47807;
    wire N__47804;
    wire N__47801;
    wire N__47796;
    wire N__47787;
    wire N__47784;
    wire N__47783;
    wire N__47782;
    wire N__47779;
    wire N__47776;
    wire N__47773;
    wire N__47770;
    wire N__47767;
    wire N__47766;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47754;
    wire N__47751;
    wire N__47742;
    wire N__47739;
    wire N__47736;
    wire N__47735;
    wire N__47732;
    wire N__47729;
    wire N__47728;
    wire N__47723;
    wire N__47720;
    wire N__47715;
    wire N__47712;
    wire N__47709;
    wire N__47706;
    wire N__47703;
    wire N__47702;
    wire N__47701;
    wire N__47700;
    wire N__47699;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47691;
    wire N__47690;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47677;
    wire N__47672;
    wire N__47669;
    wire N__47668;
    wire N__47663;
    wire N__47662;
    wire N__47659;
    wire N__47656;
    wire N__47653;
    wire N__47650;
    wire N__47645;
    wire N__47644;
    wire N__47641;
    wire N__47638;
    wire N__47635;
    wire N__47634;
    wire N__47633;
    wire N__47632;
    wire N__47631;
    wire N__47630;
    wire N__47627;
    wire N__47626;
    wire N__47619;
    wire N__47616;
    wire N__47615;
    wire N__47612;
    wire N__47611;
    wire N__47610;
    wire N__47605;
    wire N__47602;
    wire N__47597;
    wire N__47590;
    wire N__47587;
    wire N__47584;
    wire N__47579;
    wire N__47576;
    wire N__47569;
    wire N__47566;
    wire N__47559;
    wire N__47544;
    wire N__47541;
    wire N__47538;
    wire N__47537;
    wire N__47534;
    wire N__47531;
    wire N__47528;
    wire N__47527;
    wire N__47524;
    wire N__47521;
    wire N__47520;
    wire N__47517;
    wire N__47512;
    wire N__47509;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47481;
    wire N__47478;
    wire N__47477;
    wire N__47476;
    wire N__47473;
    wire N__47470;
    wire N__47467;
    wire N__47460;
    wire N__47457;
    wire N__47454;
    wire N__47453;
    wire N__47452;
    wire N__47449;
    wire N__47446;
    wire N__47443;
    wire N__47436;
    wire N__47433;
    wire N__47430;
    wire N__47429;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47419;
    wire N__47412;
    wire N__47409;
    wire N__47406;
    wire N__47405;
    wire N__47404;
    wire N__47401;
    wire N__47398;
    wire N__47395;
    wire N__47388;
    wire N__47385;
    wire N__47382;
    wire N__47381;
    wire N__47380;
    wire N__47377;
    wire N__47374;
    wire N__47371;
    wire N__47364;
    wire N__47361;
    wire N__47358;
    wire N__47357;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47347;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47333;
    wire N__47332;
    wire N__47329;
    wire N__47326;
    wire N__47323;
    wire N__47316;
    wire N__47313;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47294;
    wire N__47293;
    wire N__47290;
    wire N__47287;
    wire N__47284;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47270;
    wire N__47269;
    wire N__47266;
    wire N__47263;
    wire N__47260;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47246;
    wire N__47245;
    wire N__47242;
    wire N__47239;
    wire N__47236;
    wire N__47229;
    wire N__47226;
    wire N__47223;
    wire N__47222;
    wire N__47221;
    wire N__47218;
    wire N__47215;
    wire N__47212;
    wire N__47205;
    wire N__47202;
    wire N__47199;
    wire N__47198;
    wire N__47197;
    wire N__47194;
    wire N__47191;
    wire N__47188;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47174;
    wire N__47173;
    wire N__47170;
    wire N__47167;
    wire N__47164;
    wire N__47157;
    wire N__47154;
    wire N__47151;
    wire N__47150;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47140;
    wire N__47133;
    wire N__47130;
    wire N__47127;
    wire N__47126;
    wire N__47125;
    wire N__47122;
    wire N__47119;
    wire N__47116;
    wire N__47109;
    wire N__47106;
    wire N__47103;
    wire N__47102;
    wire N__47101;
    wire N__47098;
    wire N__47095;
    wire N__47092;
    wire N__47085;
    wire N__47082;
    wire N__47079;
    wire N__47078;
    wire N__47077;
    wire N__47074;
    wire N__47071;
    wire N__47068;
    wire N__47061;
    wire N__47058;
    wire N__47055;
    wire N__47054;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47044;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47030;
    wire N__47029;
    wire N__47026;
    wire N__47023;
    wire N__47020;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47006;
    wire N__47005;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46989;
    wire N__46986;
    wire N__46983;
    wire N__46982;
    wire N__46981;
    wire N__46978;
    wire N__46975;
    wire N__46972;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46958;
    wire N__46957;
    wire N__46954;
    wire N__46951;
    wire N__46948;
    wire N__46941;
    wire N__46938;
    wire N__46935;
    wire N__46934;
    wire N__46933;
    wire N__46930;
    wire N__46927;
    wire N__46924;
    wire N__46917;
    wire N__46914;
    wire N__46911;
    wire N__46910;
    wire N__46909;
    wire N__46906;
    wire N__46903;
    wire N__46900;
    wire N__46893;
    wire N__46890;
    wire N__46887;
    wire N__46886;
    wire N__46885;
    wire N__46882;
    wire N__46879;
    wire N__46878;
    wire N__46875;
    wire N__46874;
    wire N__46869;
    wire N__46868;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46860;
    wire N__46857;
    wire N__46854;
    wire N__46851;
    wire N__46848;
    wire N__46843;
    wire N__46840;
    wire N__46827;
    wire N__46824;
    wire N__46823;
    wire N__46822;
    wire N__46821;
    wire N__46820;
    wire N__46819;
    wire N__46818;
    wire N__46817;
    wire N__46816;
    wire N__46815;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46809;
    wire N__46808;
    wire N__46807;
    wire N__46804;
    wire N__46797;
    wire N__46794;
    wire N__46791;
    wire N__46784;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46772;
    wire N__46769;
    wire N__46768;
    wire N__46767;
    wire N__46766;
    wire N__46765;
    wire N__46764;
    wire N__46761;
    wire N__46758;
    wire N__46753;
    wire N__46752;
    wire N__46751;
    wire N__46750;
    wire N__46749;
    wire N__46748;
    wire N__46745;
    wire N__46738;
    wire N__46735;
    wire N__46728;
    wire N__46727;
    wire N__46722;
    wire N__46715;
    wire N__46712;
    wire N__46709;
    wire N__46698;
    wire N__46689;
    wire N__46686;
    wire N__46671;
    wire N__46668;
    wire N__46665;
    wire N__46662;
    wire N__46659;
    wire N__46656;
    wire N__46653;
    wire N__46650;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46631;
    wire N__46630;
    wire N__46627;
    wire N__46622;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46602;
    wire N__46599;
    wire N__46596;
    wire N__46595;
    wire N__46594;
    wire N__46591;
    wire N__46588;
    wire N__46585;
    wire N__46578;
    wire N__46575;
    wire N__46572;
    wire N__46571;
    wire N__46570;
    wire N__46567;
    wire N__46564;
    wire N__46561;
    wire N__46554;
    wire N__46551;
    wire N__46548;
    wire N__46547;
    wire N__46544;
    wire N__46541;
    wire N__46538;
    wire N__46537;
    wire N__46536;
    wire N__46533;
    wire N__46530;
    wire N__46525;
    wire N__46518;
    wire N__46515;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46491;
    wire N__46488;
    wire N__46485;
    wire N__46484;
    wire N__46481;
    wire N__46480;
    wire N__46477;
    wire N__46474;
    wire N__46473;
    wire N__46472;
    wire N__46469;
    wire N__46466;
    wire N__46463;
    wire N__46460;
    wire N__46457;
    wire N__46446;
    wire N__46445;
    wire N__46442;
    wire N__46437;
    wire N__46434;
    wire N__46431;
    wire N__46428;
    wire N__46427;
    wire N__46424;
    wire N__46423;
    wire N__46422;
    wire N__46419;
    wire N__46416;
    wire N__46413;
    wire N__46410;
    wire N__46401;
    wire N__46400;
    wire N__46399;
    wire N__46396;
    wire N__46391;
    wire N__46386;
    wire N__46383;
    wire N__46382;
    wire N__46379;
    wire N__46376;
    wire N__46373;
    wire N__46368;
    wire N__46367;
    wire N__46366;
    wire N__46359;
    wire N__46356;
    wire N__46353;
    wire N__46350;
    wire N__46347;
    wire N__46346;
    wire N__46345;
    wire N__46344;
    wire N__46341;
    wire N__46338;
    wire N__46333;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46317;
    wire N__46314;
    wire N__46311;
    wire N__46310;
    wire N__46307;
    wire N__46304;
    wire N__46299;
    wire N__46298;
    wire N__46295;
    wire N__46294;
    wire N__46291;
    wire N__46284;
    wire N__46281;
    wire N__46278;
    wire N__46277;
    wire N__46274;
    wire N__46273;
    wire N__46270;
    wire N__46269;
    wire N__46266;
    wire N__46263;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46241;
    wire N__46236;
    wire N__46233;
    wire N__46232;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46206;
    wire N__46203;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46193;
    wire N__46190;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46174;
    wire N__46171;
    wire N__46166;
    wire N__46163;
    wire N__46162;
    wire N__46159;
    wire N__46156;
    wire N__46153;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46139;
    wire N__46138;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46112;
    wire N__46109;
    wire N__46106;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46096;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46068;
    wire N__46063;
    wire N__46056;
    wire N__46053;
    wire N__46052;
    wire N__46049;
    wire N__46046;
    wire N__46045;
    wire N__46042;
    wire N__46039;
    wire N__46036;
    wire N__46029;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46013;
    wire N__46012;
    wire N__46011;
    wire N__46010;
    wire N__46009;
    wire N__46008;
    wire N__46007;
    wire N__46006;
    wire N__46005;
    wire N__46004;
    wire N__46003;
    wire N__46002;
    wire N__46001;
    wire N__46000;
    wire N__45999;
    wire N__45998;
    wire N__45997;
    wire N__45996;
    wire N__45995;
    wire N__45994;
    wire N__45993;
    wire N__45992;
    wire N__45989;
    wire N__45988;
    wire N__45987;
    wire N__45986;
    wire N__45983;
    wire N__45982;
    wire N__45981;
    wire N__45980;
    wire N__45977;
    wire N__45976;
    wire N__45975;
    wire N__45974;
    wire N__45965;
    wire N__45956;
    wire N__45955;
    wire N__45954;
    wire N__45953;
    wire N__45952;
    wire N__45949;
    wire N__45948;
    wire N__45947;
    wire N__45946;
    wire N__45945;
    wire N__45944;
    wire N__45943;
    wire N__45942;
    wire N__45941;
    wire N__45940;
    wire N__45939;
    wire N__45936;
    wire N__45935;
    wire N__45932;
    wire N__45931;
    wire N__45928;
    wire N__45927;
    wire N__45924;
    wire N__45923;
    wire N__45920;
    wire N__45919;
    wire N__45916;
    wire N__45915;
    wire N__45912;
    wire N__45911;
    wire N__45910;
    wire N__45909;
    wire N__45908;
    wire N__45907;
    wire N__45906;
    wire N__45905;
    wire N__45904;
    wire N__45903;
    wire N__45902;
    wire N__45901;
    wire N__45900;
    wire N__45897;
    wire N__45896;
    wire N__45893;
    wire N__45892;
    wire N__45889;
    wire N__45888;
    wire N__45887;
    wire N__45886;
    wire N__45885;
    wire N__45884;
    wire N__45883;
    wire N__45882;
    wire N__45877;
    wire N__45876;
    wire N__45875;
    wire N__45874;
    wire N__45871;
    wire N__45864;
    wire N__45853;
    wire N__45852;
    wire N__45849;
    wire N__45848;
    wire N__45845;
    wire N__45844;
    wire N__45843;
    wire N__45842;
    wire N__45841;
    wire N__45840;
    wire N__45835;
    wire N__45822;
    wire N__45811;
    wire N__45806;
    wire N__45805;
    wire N__45804;
    wire N__45803;
    wire N__45802;
    wire N__45801;
    wire N__45784;
    wire N__45767;
    wire N__45764;
    wire N__45763;
    wire N__45760;
    wire N__45759;
    wire N__45756;
    wire N__45755;
    wire N__45752;
    wire N__45751;
    wire N__45750;
    wire N__45749;
    wire N__45748;
    wire N__45747;
    wire N__45744;
    wire N__45743;
    wire N__45740;
    wire N__45739;
    wire N__45736;
    wire N__45735;
    wire N__45732;
    wire N__45731;
    wire N__45728;
    wire N__45727;
    wire N__45724;
    wire N__45723;
    wire N__45720;
    wire N__45719;
    wire N__45706;
    wire N__45697;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45685;
    wire N__45682;
    wire N__45681;
    wire N__45680;
    wire N__45679;
    wire N__45676;
    wire N__45675;
    wire N__45674;
    wire N__45673;
    wire N__45672;
    wire N__45667;
    wire N__45664;
    wire N__45653;
    wire N__45650;
    wire N__45649;
    wire N__45646;
    wire N__45645;
    wire N__45642;
    wire N__45641;
    wire N__45638;
    wire N__45637;
    wire N__45628;
    wire N__45617;
    wire N__45612;
    wire N__45595;
    wire N__45592;
    wire N__45591;
    wire N__45588;
    wire N__45587;
    wire N__45584;
    wire N__45583;
    wire N__45568;
    wire N__45551;
    wire N__45548;
    wire N__45543;
    wire N__45538;
    wire N__45523;
    wire N__45516;
    wire N__45509;
    wire N__45492;
    wire N__45483;
    wire N__45470;
    wire N__45463;
    wire N__45444;
    wire N__45443;
    wire N__45442;
    wire N__45441;
    wire N__45440;
    wire N__45439;
    wire N__45438;
    wire N__45437;
    wire N__45436;
    wire N__45435;
    wire N__45434;
    wire N__45433;
    wire N__45432;
    wire N__45431;
    wire N__45430;
    wire N__45429;
    wire N__45428;
    wire N__45427;
    wire N__45426;
    wire N__45425;
    wire N__45424;
    wire N__45423;
    wire N__45422;
    wire N__45421;
    wire N__45420;
    wire N__45419;
    wire N__45418;
    wire N__45417;
    wire N__45416;
    wire N__45415;
    wire N__45414;
    wire N__45413;
    wire N__45412;
    wire N__45411;
    wire N__45410;
    wire N__45409;
    wire N__45408;
    wire N__45407;
    wire N__45406;
    wire N__45405;
    wire N__45404;
    wire N__45403;
    wire N__45400;
    wire N__45399;
    wire N__45398;
    wire N__45397;
    wire N__45396;
    wire N__45395;
    wire N__45394;
    wire N__45393;
    wire N__45392;
    wire N__45389;
    wire N__45378;
    wire N__45365;
    wire N__45364;
    wire N__45355;
    wire N__45346;
    wire N__45345;
    wire N__45344;
    wire N__45343;
    wire N__45342;
    wire N__45341;
    wire N__45340;
    wire N__45339;
    wire N__45338;
    wire N__45333;
    wire N__45324;
    wire N__45313;
    wire N__45306;
    wire N__45303;
    wire N__45302;
    wire N__45301;
    wire N__45300;
    wire N__45299;
    wire N__45298;
    wire N__45297;
    wire N__45286;
    wire N__45283;
    wire N__45268;
    wire N__45267;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45257;
    wire N__45252;
    wire N__45251;
    wire N__45250;
    wire N__45249;
    wire N__45246;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45221;
    wire N__45216;
    wire N__45213;
    wire N__45208;
    wire N__45195;
    wire N__45192;
    wire N__45187;
    wire N__45182;
    wire N__45173;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45145;
    wire N__45126;
    wire N__45123;
    wire N__45122;
    wire N__45119;
    wire N__45116;
    wire N__45115;
    wire N__45112;
    wire N__45107;
    wire N__45102;
    wire N__45101;
    wire N__45096;
    wire N__45095;
    wire N__45094;
    wire N__45091;
    wire N__45086;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45057;
    wire N__45054;
    wire N__45051;
    wire N__45048;
    wire N__45045;
    wire N__45042;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45032;
    wire N__45029;
    wire N__45026;
    wire N__45021;
    wire N__45018;
    wire N__45015;
    wire N__45012;
    wire N__45009;
    wire N__45006;
    wire N__45003;
    wire N__45002;
    wire N__44999;
    wire N__44998;
    wire N__44995;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44982;
    wire N__44977;
    wire N__44974;
    wire N__44969;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44957;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44924;
    wire N__44921;
    wire N__44918;
    wire N__44917;
    wire N__44912;
    wire N__44909;
    wire N__44906;
    wire N__44901;
    wire N__44900;
    wire N__44899;
    wire N__44898;
    wire N__44893;
    wire N__44890;
    wire N__44887;
    wire N__44884;
    wire N__44881;
    wire N__44878;
    wire N__44875;
    wire N__44872;
    wire N__44869;
    wire N__44862;
    wire N__44859;
    wire N__44858;
    wire N__44857;
    wire N__44852;
    wire N__44849;
    wire N__44846;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44825;
    wire N__44822;
    wire N__44819;
    wire N__44816;
    wire N__44813;
    wire N__44812;
    wire N__44809;
    wire N__44806;
    wire N__44803;
    wire N__44802;
    wire N__44797;
    wire N__44792;
    wire N__44789;
    wire N__44786;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44774;
    wire N__44773;
    wire N__44770;
    wire N__44767;
    wire N__44764;
    wire N__44757;
    wire N__44754;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44741;
    wire N__44740;
    wire N__44737;
    wire N__44734;
    wire N__44733;
    wire N__44732;
    wire N__44729;
    wire N__44726;
    wire N__44723;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44706;
    wire N__44701;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44676;
    wire N__44675;
    wire N__44672;
    wire N__44671;
    wire N__44668;
    wire N__44665;
    wire N__44662;
    wire N__44659;
    wire N__44656;
    wire N__44653;
    wire N__44652;
    wire N__44649;
    wire N__44644;
    wire N__44641;
    wire N__44634;
    wire N__44631;
    wire N__44628;
    wire N__44627;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44617;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44601;
    wire N__44598;
    wire N__44597;
    wire N__44596;
    wire N__44595;
    wire N__44594;
    wire N__44593;
    wire N__44592;
    wire N__44591;
    wire N__44590;
    wire N__44589;
    wire N__44588;
    wire N__44587;
    wire N__44586;
    wire N__44585;
    wire N__44584;
    wire N__44583;
    wire N__44582;
    wire N__44581;
    wire N__44580;
    wire N__44577;
    wire N__44576;
    wire N__44575;
    wire N__44574;
    wire N__44571;
    wire N__44570;
    wire N__44569;
    wire N__44566;
    wire N__44565;
    wire N__44560;
    wire N__44559;
    wire N__44556;
    wire N__44555;
    wire N__44554;
    wire N__44551;
    wire N__44548;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44535;
    wire N__44532;
    wire N__44531;
    wire N__44528;
    wire N__44525;
    wire N__44524;
    wire N__44523;
    wire N__44522;
    wire N__44519;
    wire N__44518;
    wire N__44517;
    wire N__44516;
    wire N__44515;
    wire N__44514;
    wire N__44513;
    wire N__44512;
    wire N__44511;
    wire N__44510;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44496;
    wire N__44495;
    wire N__44492;
    wire N__44481;
    wire N__44478;
    wire N__44475;
    wire N__44474;
    wire N__44461;
    wire N__44458;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44444;
    wire N__44427;
    wire N__44420;
    wire N__44417;
    wire N__44414;
    wire N__44407;
    wire N__44404;
    wire N__44401;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44386;
    wire N__44381;
    wire N__44380;
    wire N__44377;
    wire N__44376;
    wire N__44375;
    wire N__44374;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44358;
    wire N__44353;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44325;
    wire N__44314;
    wire N__44305;
    wire N__44300;
    wire N__44283;
    wire N__44282;
    wire N__44279;
    wire N__44276;
    wire N__44273;
    wire N__44270;
    wire N__44269;
    wire N__44266;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44247;
    wire N__44244;
    wire N__44243;
    wire N__44240;
    wire N__44237;
    wire N__44236;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44220;
    wire N__44217;
    wire N__44216;
    wire N__44213;
    wire N__44212;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44199;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44159;
    wire N__44156;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44143;
    wire N__44136;
    wire N__44135;
    wire N__44134;
    wire N__44133;
    wire N__44132;
    wire N__44131;
    wire N__44130;
    wire N__44129;
    wire N__44128;
    wire N__44109;
    wire N__44106;
    wire N__44103;
    wire N__44102;
    wire N__44099;
    wire N__44094;
    wire N__44093;
    wire N__44090;
    wire N__44087;
    wire N__44086;
    wire N__44081;
    wire N__44078;
    wire N__44075;
    wire N__44070;
    wire N__44067;
    wire N__44064;
    wire N__44061;
    wire N__44058;
    wire N__44055;
    wire N__44054;
    wire N__44053;
    wire N__44052;
    wire N__44051;
    wire N__44050;
    wire N__44049;
    wire N__44048;
    wire N__44047;
    wire N__44046;
    wire N__44045;
    wire N__44042;
    wire N__44041;
    wire N__44040;
    wire N__44039;
    wire N__44038;
    wire N__44037;
    wire N__44036;
    wire N__44033;
    wire N__44028;
    wire N__44025;
    wire N__44024;
    wire N__44023;
    wire N__44022;
    wire N__44021;
    wire N__44020;
    wire N__44019;
    wire N__44018;
    wire N__44017;
    wire N__44004;
    wire N__44001;
    wire N__43992;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43975;
    wire N__43960;
    wire N__43955;
    wire N__43952;
    wire N__43945;
    wire N__43932;
    wire N__43931;
    wire N__43928;
    wire N__43927;
    wire N__43920;
    wire N__43917;
    wire N__43916;
    wire N__43915;
    wire N__43914;
    wire N__43907;
    wire N__43904;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43860;
    wire N__43857;
    wire N__43854;
    wire N__43851;
    wire N__43850;
    wire N__43847;
    wire N__43844;
    wire N__43843;
    wire N__43842;
    wire N__43841;
    wire N__43836;
    wire N__43831;
    wire N__43828;
    wire N__43823;
    wire N__43818;
    wire N__43817;
    wire N__43816;
    wire N__43813;
    wire N__43808;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43794;
    wire N__43791;
    wire N__43788;
    wire N__43785;
    wire N__43782;
    wire N__43779;
    wire N__43776;
    wire N__43775;
    wire N__43774;
    wire N__43773;
    wire N__43770;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43750;
    wire N__43747;
    wire N__43740;
    wire N__43737;
    wire N__43736;
    wire N__43733;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43718;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43674;
    wire N__43671;
    wire N__43668;
    wire N__43663;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43647;
    wire N__43646;
    wire N__43643;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43608;
    wire N__43607;
    wire N__43604;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43580;
    wire N__43579;
    wire N__43576;
    wire N__43573;
    wire N__43570;
    wire N__43563;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43553;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43536;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43489;
    wire N__43488;
    wire N__43485;
    wire N__43482;
    wire N__43477;
    wire N__43474;
    wire N__43469;
    wire N__43464;
    wire N__43461;
    wire N__43458;
    wire N__43457;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43440;
    wire N__43437;
    wire N__43434;
    wire N__43431;
    wire N__43428;
    wire N__43425;
    wire N__43422;
    wire N__43421;
    wire N__43418;
    wire N__43415;
    wire N__43414;
    wire N__43413;
    wire N__43410;
    wire N__43407;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43393;
    wire N__43386;
    wire N__43385;
    wire N__43382;
    wire N__43379;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43364;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43335;
    wire N__43334;
    wire N__43331;
    wire N__43328;
    wire N__43327;
    wire N__43322;
    wire N__43319;
    wire N__43314;
    wire N__43313;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43302;
    wire N__43299;
    wire N__43296;
    wire N__43291;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43272;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43241;
    wire N__43238;
    wire N__43235;
    wire N__43230;
    wire N__43227;
    wire N__43224;
    wire N__43221;
    wire N__43220;
    wire N__43217;
    wire N__43214;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43187;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43169;
    wire N__43166;
    wire N__43163;
    wire N__43158;
    wire N__43155;
    wire N__43152;
    wire N__43151;
    wire N__43148;
    wire N__43145;
    wire N__43142;
    wire N__43139;
    wire N__43134;
    wire N__43131;
    wire N__43128;
    wire N__43125;
    wire N__43124;
    wire N__43121;
    wire N__43118;
    wire N__43113;
    wire N__43110;
    wire N__43109;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43092;
    wire N__43089;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43071;
    wire N__43068;
    wire N__43067;
    wire N__43066;
    wire N__43063;
    wire N__43062;
    wire N__43057;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43041;
    wire N__43038;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43025;
    wire N__43024;
    wire N__43019;
    wire N__43016;
    wire N__43011;
    wire N__43008;
    wire N__43007;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42981;
    wire N__42978;
    wire N__42975;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42967;
    wire N__42964;
    wire N__42961;
    wire N__42958;
    wire N__42951;
    wire N__42948;
    wire N__42945;
    wire N__42942;
    wire N__42941;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42924;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42908;
    wire N__42905;
    wire N__42902;
    wire N__42897;
    wire N__42894;
    wire N__42891;
    wire N__42890;
    wire N__42889;
    wire N__42886;
    wire N__42881;
    wire N__42876;
    wire N__42873;
    wire N__42870;
    wire N__42869;
    wire N__42868;
    wire N__42865;
    wire N__42860;
    wire N__42857;
    wire N__42854;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42831;
    wire N__42830;
    wire N__42829;
    wire N__42826;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42807;
    wire N__42798;
    wire N__42795;
    wire N__42792;
    wire N__42791;
    wire N__42788;
    wire N__42785;
    wire N__42780;
    wire N__42777;
    wire N__42774;
    wire N__42773;
    wire N__42770;
    wire N__42767;
    wire N__42762;
    wire N__42759;
    wire N__42756;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42743;
    wire N__42738;
    wire N__42735;
    wire N__42732;
    wire N__42729;
    wire N__42728;
    wire N__42725;
    wire N__42722;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42696;
    wire N__42693;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42671;
    wire N__42668;
    wire N__42665;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42653;
    wire N__42652;
    wire N__42649;
    wire N__42644;
    wire N__42639;
    wire N__42636;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42617;
    wire N__42614;
    wire N__42611;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42599;
    wire N__42596;
    wire N__42593;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42578;
    wire N__42575;
    wire N__42572;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42560;
    wire N__42557;
    wire N__42556;
    wire N__42555;
    wire N__42554;
    wire N__42551;
    wire N__42548;
    wire N__42545;
    wire N__42542;
    wire N__42539;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42521;
    wire N__42518;
    wire N__42517;
    wire N__42516;
    wire N__42515;
    wire N__42512;
    wire N__42509;
    wire N__42506;
    wire N__42503;
    wire N__42500;
    wire N__42489;
    wire N__42486;
    wire N__42485;
    wire N__42482;
    wire N__42479;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42467;
    wire N__42464;
    wire N__42461;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42449;
    wire N__42446;
    wire N__42443;
    wire N__42442;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42430;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42404;
    wire N__42401;
    wire N__42398;
    wire N__42397;
    wire N__42392;
    wire N__42389;
    wire N__42388;
    wire N__42385;
    wire N__42382;
    wire N__42379;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42356;
    wire N__42353;
    wire N__42350;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42335;
    wire N__42334;
    wire N__42331;
    wire N__42328;
    wire N__42325;
    wire N__42322;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42276;
    wire N__42273;
    wire N__42270;
    wire N__42267;
    wire N__42266;
    wire N__42263;
    wire N__42260;
    wire N__42257;
    wire N__42254;
    wire N__42253;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42239;
    wire N__42234;
    wire N__42231;
    wire N__42230;
    wire N__42229;
    wire N__42226;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42213;
    wire N__42204;
    wire N__42203;
    wire N__42200;
    wire N__42199;
    wire N__42196;
    wire N__42193;
    wire N__42190;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42174;
    wire N__42171;
    wire N__42170;
    wire N__42169;
    wire N__42168;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42158;
    wire N__42155;
    wire N__42152;
    wire N__42149;
    wire N__42146;
    wire N__42143;
    wire N__42132;
    wire N__42129;
    wire N__42128;
    wire N__42127;
    wire N__42124;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42106;
    wire N__42105;
    wire N__42102;
    wire N__42097;
    wire N__42094;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42048;
    wire N__42045;
    wire N__42042;
    wire N__42039;
    wire N__42036;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41991;
    wire N__41988;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41919;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41859;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41841;
    wire N__41838;
    wire N__41835;
    wire N__41832;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41787;
    wire N__41784;
    wire N__41781;
    wire N__41780;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41765;
    wire N__41762;
    wire N__41761;
    wire N__41756;
    wire N__41753;
    wire N__41752;
    wire N__41749;
    wire N__41744;
    wire N__41739;
    wire N__41736;
    wire N__41735;
    wire N__41734;
    wire N__41731;
    wire N__41728;
    wire N__41725;
    wire N__41720;
    wire N__41717;
    wire N__41714;
    wire N__41709;
    wire N__41708;
    wire N__41705;
    wire N__41702;
    wire N__41701;
    wire N__41698;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41680;
    wire N__41677;
    wire N__41674;
    wire N__41671;
    wire N__41666;
    wire N__41661;
    wire N__41658;
    wire N__41657;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41642;
    wire N__41637;
    wire N__41634;
    wire N__41633;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41616;
    wire N__41613;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41600;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41577;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41556;
    wire N__41553;
    wire N__41550;
    wire N__41549;
    wire N__41548;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41499;
    wire N__41496;
    wire N__41493;
    wire N__41490;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41480;
    wire N__41477;
    wire N__41474;
    wire N__41473;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41459;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41414;
    wire N__41409;
    wire N__41406;
    wire N__41403;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41383;
    wire N__41380;
    wire N__41375;
    wire N__41370;
    wire N__41367;
    wire N__41364;
    wire N__41361;
    wire N__41358;
    wire N__41357;
    wire N__41356;
    wire N__41349;
    wire N__41346;
    wire N__41343;
    wire N__41340;
    wire N__41337;
    wire N__41334;
    wire N__41331;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41280;
    wire N__41277;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41252;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41204;
    wire N__41203;
    wire N__41200;
    wire N__41197;
    wire N__41194;
    wire N__41189;
    wire N__41184;
    wire N__41181;
    wire N__41178;
    wire N__41175;
    wire N__41172;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41149;
    wire N__41146;
    wire N__41141;
    wire N__41138;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41102;
    wire N__41099;
    wire N__41096;
    wire N__41093;
    wire N__41090;
    wire N__41089;
    wire N__41088;
    wire N__41085;
    wire N__41082;
    wire N__41077;
    wire N__41074;
    wire N__41069;
    wire N__41064;
    wire N__41063;
    wire N__41060;
    wire N__41057;
    wire N__41056;
    wire N__41053;
    wire N__41050;
    wire N__41049;
    wire N__41046;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41018;
    wire N__41013;
    wire N__41010;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__40998;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40986;
    wire N__40983;
    wire N__40980;
    wire N__40979;
    wire N__40978;
    wire N__40975;
    wire N__40972;
    wire N__40969;
    wire N__40962;
    wire N__40959;
    wire N__40956;
    wire N__40953;
    wire N__40950;
    wire N__40947;
    wire N__40944;
    wire N__40943;
    wire N__40942;
    wire N__40939;
    wire N__40934;
    wire N__40931;
    wire N__40926;
    wire N__40923;
    wire N__40922;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40914;
    wire N__40911;
    wire N__40908;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40893;
    wire N__40884;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40868;
    wire N__40867;
    wire N__40866;
    wire N__40865;
    wire N__40864;
    wire N__40861;
    wire N__40860;
    wire N__40859;
    wire N__40858;
    wire N__40855;
    wire N__40850;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40838;
    wire N__40835;
    wire N__40832;
    wire N__40831;
    wire N__40828;
    wire N__40825;
    wire N__40820;
    wire N__40815;
    wire N__40812;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40798;
    wire N__40785;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40775;
    wire N__40770;
    wire N__40767;
    wire N__40766;
    wire N__40763;
    wire N__40760;
    wire N__40757;
    wire N__40754;
    wire N__40751;
    wire N__40746;
    wire N__40745;
    wire N__40742;
    wire N__40739;
    wire N__40734;
    wire N__40733;
    wire N__40730;
    wire N__40727;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40707;
    wire N__40704;
    wire N__40703;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40681;
    wire N__40678;
    wire N__40673;
    wire N__40668;
    wire N__40667;
    wire N__40666;
    wire N__40661;
    wire N__40658;
    wire N__40655;
    wire N__40652;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40635;
    wire N__40632;
    wire N__40631;
    wire N__40628;
    wire N__40625;
    wire N__40620;
    wire N__40617;
    wire N__40616;
    wire N__40613;
    wire N__40610;
    wire N__40605;
    wire N__40604;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40586;
    wire N__40583;
    wire N__40580;
    wire N__40577;
    wire N__40574;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40560;
    wire N__40559;
    wire N__40556;
    wire N__40553;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40538;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40521;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40509;
    wire N__40506;
    wire N__40505;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40493;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40481;
    wire N__40476;
    wire N__40473;
    wire N__40470;
    wire N__40469;
    wire N__40466;
    wire N__40463;
    wire N__40458;
    wire N__40455;
    wire N__40452;
    wire N__40449;
    wire N__40446;
    wire N__40445;
    wire N__40442;
    wire N__40439;
    wire N__40434;
    wire N__40433;
    wire N__40430;
    wire N__40427;
    wire N__40424;
    wire N__40419;
    wire N__40416;
    wire N__40415;
    wire N__40414;
    wire N__40411;
    wire N__40408;
    wire N__40405;
    wire N__40398;
    wire N__40397;
    wire N__40394;
    wire N__40391;
    wire N__40386;
    wire N__40383;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40319;
    wire N__40318;
    wire N__40315;
    wire N__40314;
    wire N__40311;
    wire N__40308;
    wire N__40305;
    wire N__40302;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40278;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40245;
    wire N__40244;
    wire N__40243;
    wire N__40240;
    wire N__40235;
    wire N__40230;
    wire N__40227;
    wire N__40224;
    wire N__40223;
    wire N__40222;
    wire N__40219;
    wire N__40216;
    wire N__40213;
    wire N__40208;
    wire N__40205;
    wire N__40204;
    wire N__40201;
    wire N__40198;
    wire N__40195;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40152;
    wire N__40149;
    wire N__40146;
    wire N__40143;
    wire N__40140;
    wire N__40137;
    wire N__40134;
    wire N__40131;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40123;
    wire N__40120;
    wire N__40117;
    wire N__40114;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40092;
    wire N__40089;
    wire N__40086;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40074;
    wire N__40073;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40062;
    wire N__40059;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40049;
    wire N__40046;
    wire N__40043;
    wire N__40040;
    wire N__40035;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__40002;
    wire N__39999;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39980;
    wire N__39977;
    wire N__39974;
    wire N__39973;
    wire N__39968;
    wire N__39965;
    wire N__39960;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39947;
    wire N__39942;
    wire N__39941;
    wire N__39940;
    wire N__39937;
    wire N__39932;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39863;
    wire N__39860;
    wire N__39859;
    wire N__39852;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39806;
    wire N__39803;
    wire N__39802;
    wire N__39795;
    wire N__39792;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39759;
    wire N__39756;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39744;
    wire N__39741;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39729;
    wire N__39726;
    wire N__39723;
    wire N__39720;
    wire N__39717;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39683;
    wire N__39682;
    wire N__39681;
    wire N__39678;
    wire N__39673;
    wire N__39668;
    wire N__39665;
    wire N__39662;
    wire N__39659;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39636;
    wire N__39633;
    wire N__39630;
    wire N__39627;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39612;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39600;
    wire N__39599;
    wire N__39596;
    wire N__39593;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39578;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39561;
    wire N__39560;
    wire N__39559;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39534;
    wire N__39531;
    wire N__39528;
    wire N__39525;
    wire N__39524;
    wire N__39523;
    wire N__39520;
    wire N__39515;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39498;
    wire N__39495;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39425;
    wire N__39424;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39408;
    wire N__39407;
    wire N__39406;
    wire N__39403;
    wire N__39398;
    wire N__39393;
    wire N__39390;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39374;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39359;
    wire N__39358;
    wire N__39355;
    wire N__39354;
    wire N__39351;
    wire N__39348;
    wire N__39345;
    wire N__39342;
    wire N__39339;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39323;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39313;
    wire N__39310;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39290;
    wire N__39287;
    wire N__39284;
    wire N__39279;
    wire N__39278;
    wire N__39275;
    wire N__39272;
    wire N__39267;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39167;
    wire N__39164;
    wire N__39161;
    wire N__39158;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39123;
    wire N__39120;
    wire N__39117;
    wire N__39116;
    wire N__39113;
    wire N__39110;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39090;
    wire N__39089;
    wire N__39086;
    wire N__39083;
    wire N__39078;
    wire N__39075;
    wire N__39072;
    wire N__39069;
    wire N__39068;
    wire N__39065;
    wire N__39062;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39045;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39021;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39000;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38978;
    wire N__38975;
    wire N__38972;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38957;
    wire N__38954;
    wire N__38951;
    wire N__38948;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38921;
    wire N__38918;
    wire N__38915;
    wire N__38910;
    wire N__38907;
    wire N__38904;
    wire N__38901;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38889;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38879;
    wire N__38876;
    wire N__38873;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38858;
    wire N__38855;
    wire N__38852;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38813;
    wire N__38812;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38796;
    wire N__38793;
    wire N__38792;
    wire N__38787;
    wire N__38784;
    wire N__38783;
    wire N__38782;
    wire N__38779;
    wire N__38774;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38724;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38672;
    wire N__38669;
    wire N__38666;
    wire N__38661;
    wire N__38660;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38648;
    wire N__38643;
    wire N__38642;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38609;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38521;
    wire N__38520;
    wire N__38519;
    wire N__38518;
    wire N__38515;
    wire N__38514;
    wire N__38513;
    wire N__38512;
    wire N__38509;
    wire N__38500;
    wire N__38499;
    wire N__38498;
    wire N__38497;
    wire N__38496;
    wire N__38495;
    wire N__38494;
    wire N__38491;
    wire N__38484;
    wire N__38479;
    wire N__38468;
    wire N__38465;
    wire N__38454;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38337;
    wire N__38334;
    wire N__38331;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38282;
    wire N__38281;
    wire N__38280;
    wire N__38279;
    wire N__38278;
    wire N__38277;
    wire N__38276;
    wire N__38275;
    wire N__38274;
    wire N__38271;
    wire N__38270;
    wire N__38267;
    wire N__38260;
    wire N__38251;
    wire N__38250;
    wire N__38249;
    wire N__38248;
    wire N__38247;
    wire N__38246;
    wire N__38245;
    wire N__38244;
    wire N__38243;
    wire N__38240;
    wire N__38237;
    wire N__38236;
    wire N__38233;
    wire N__38226;
    wire N__38223;
    wire N__38216;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38200;
    wire N__38199;
    wire N__38198;
    wire N__38195;
    wire N__38194;
    wire N__38193;
    wire N__38192;
    wire N__38189;
    wire N__38180;
    wire N__38175;
    wire N__38172;
    wire N__38167;
    wire N__38164;
    wire N__38163;
    wire N__38162;
    wire N__38161;
    wire N__38158;
    wire N__38157;
    wire N__38154;
    wire N__38153;
    wire N__38150;
    wire N__38149;
    wire N__38148;
    wire N__38147;
    wire N__38146;
    wire N__38145;
    wire N__38144;
    wire N__38143;
    wire N__38142;
    wire N__38141;
    wire N__38140;
    wire N__38139;
    wire N__38138;
    wire N__38135;
    wire N__38132;
    wire N__38125;
    wire N__38122;
    wire N__38117;
    wire N__38102;
    wire N__38099;
    wire N__38098;
    wire N__38095;
    wire N__38094;
    wire N__38091;
    wire N__38090;
    wire N__38087;
    wire N__38086;
    wire N__38083;
    wire N__38082;
    wire N__38079;
    wire N__38078;
    wire N__38075;
    wire N__38074;
    wire N__38071;
    wire N__38070;
    wire N__38069;
    wire N__38066;
    wire N__38065;
    wire N__38062;
    wire N__38061;
    wire N__38058;
    wire N__38057;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38043;
    wire N__38040;
    wire N__38023;
    wire N__38006;
    wire N__37991;
    wire N__37986;
    wire N__37981;
    wire N__37972;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37915;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37899;
    wire N__37896;
    wire N__37895;
    wire N__37892;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37881;
    wire N__37878;
    wire N__37877;
    wire N__37874;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37855;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37821;
    wire N__37818;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37755;
    wire N__37752;
    wire N__37751;
    wire N__37748;
    wire N__37745;
    wire N__37740;
    wire N__37737;
    wire N__37736;
    wire N__37733;
    wire N__37730;
    wire N__37727;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37701;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37671;
    wire N__37668;
    wire N__37667;
    wire N__37662;
    wire N__37659;
    wire N__37656;
    wire N__37655;
    wire N__37654;
    wire N__37653;
    wire N__37652;
    wire N__37649;
    wire N__37644;
    wire N__37639;
    wire N__37632;
    wire N__37631;
    wire N__37630;
    wire N__37627;
    wire N__37626;
    wire N__37625;
    wire N__37622;
    wire N__37613;
    wire N__37608;
    wire N__37607;
    wire N__37604;
    wire N__37601;
    wire N__37596;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37581;
    wire N__37578;
    wire N__37575;
    wire N__37572;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37546;
    wire N__37545;
    wire N__37540;
    wire N__37535;
    wire N__37532;
    wire N__37527;
    wire N__37524;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37498;
    wire N__37491;
    wire N__37488;
    wire N__37485;
    wire N__37484;
    wire N__37483;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37470;
    wire N__37467;
    wire N__37458;
    wire N__37457;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37444;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37413;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37383;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37341;
    wire N__37338;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37245;
    wire N__37242;
    wire N__37239;
    wire N__37236;
    wire N__37235;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37221;
    wire N__37218;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37203;
    wire N__37200;
    wire N__37199;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37185;
    wire N__37182;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37158;
    wire N__37155;
    wire N__37152;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37137;
    wire N__37134;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37119;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37104;
    wire N__37101;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37086;
    wire N__37083;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37068;
    wire N__37065;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37055;
    wire N__37050;
    wire N__37047;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37032;
    wire N__37029;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36993;
    wire N__36990;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36975;
    wire N__36972;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36930;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36914;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36897;
    wire N__36894;
    wire N__36891;
    wire N__36888;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36873;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36836;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36818;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36792;
    wire N__36791;
    wire N__36788;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36768;
    wire N__36765;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36730;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36714;
    wire N__36711;
    wire N__36710;
    wire N__36709;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36693;
    wire N__36690;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36680;
    wire N__36675;
    wire N__36672;
    wire N__36671;
    wire N__36670;
    wire N__36669;
    wire N__36668;
    wire N__36667;
    wire N__36666;
    wire N__36665;
    wire N__36664;
    wire N__36663;
    wire N__36658;
    wire N__36657;
    wire N__36656;
    wire N__36655;
    wire N__36654;
    wire N__36653;
    wire N__36652;
    wire N__36651;
    wire N__36650;
    wire N__36649;
    wire N__36648;
    wire N__36647;
    wire N__36646;
    wire N__36637;
    wire N__36636;
    wire N__36635;
    wire N__36634;
    wire N__36633;
    wire N__36632;
    wire N__36631;
    wire N__36630;
    wire N__36629;
    wire N__36620;
    wire N__36617;
    wire N__36608;
    wire N__36599;
    wire N__36590;
    wire N__36587;
    wire N__36578;
    wire N__36569;
    wire N__36558;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36528;
    wire N__36525;
    wire N__36524;
    wire N__36523;
    wire N__36520;
    wire N__36517;
    wire N__36516;
    wire N__36513;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36497;
    wire N__36494;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36474;
    wire N__36473;
    wire N__36470;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36460;
    wire N__36453;
    wire N__36450;
    wire N__36449;
    wire N__36444;
    wire N__36443;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36429;
    wire N__36426;
    wire N__36425;
    wire N__36424;
    wire N__36419;
    wire N__36416;
    wire N__36413;
    wire N__36408;
    wire N__36405;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36393;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36378;
    wire N__36375;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36367;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36351;
    wire N__36348;
    wire N__36347;
    wire N__36346;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36330;
    wire N__36327;
    wire N__36326;
    wire N__36323;
    wire N__36320;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36305;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36293;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36261;
    wire N__36260;
    wire N__36257;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36240;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36230;
    wire N__36227;
    wire N__36226;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36210;
    wire N__36207;
    wire N__36206;
    wire N__36201;
    wire N__36200;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36186;
    wire N__36183;
    wire N__36182;
    wire N__36181;
    wire N__36176;
    wire N__36173;
    wire N__36170;
    wire N__36165;
    wire N__36162;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36150;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36140;
    wire N__36135;
    wire N__36132;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36124;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36108;
    wire N__36105;
    wire N__36104;
    wire N__36103;
    wire N__36098;
    wire N__36095;
    wire N__36092;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36073;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36050;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36013;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35990;
    wire N__35987;
    wire N__35986;
    wire N__35983;
    wire N__35980;
    wire N__35977;
    wire N__35974;
    wire N__35971;
    wire N__35964;
    wire N__35961;
    wire N__35960;
    wire N__35959;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35943;
    wire N__35940;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35932;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35916;
    wire N__35913;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35901;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35886;
    wire N__35883;
    wire N__35882;
    wire N__35879;
    wire N__35876;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35861;
    wire N__35856;
    wire N__35853;
    wire N__35850;
    wire N__35849;
    wire N__35846;
    wire N__35845;
    wire N__35842;
    wire N__35839;
    wire N__35836;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35813;
    wire N__35810;
    wire N__35807;
    wire N__35806;
    wire N__35801;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35784;
    wire N__35781;
    wire N__35780;
    wire N__35779;
    wire N__35776;
    wire N__35775;
    wire N__35770;
    wire N__35767;
    wire N__35764;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35750;
    wire N__35749;
    wire N__35748;
    wire N__35745;
    wire N__35740;
    wire N__35737;
    wire N__35734;
    wire N__35727;
    wire N__35724;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35700;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35679;
    wire N__35678;
    wire N__35673;
    wire N__35670;
    wire N__35669;
    wire N__35668;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35652;
    wire N__35651;
    wire N__35650;
    wire N__35649;
    wire N__35646;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35636;
    wire N__35633;
    wire N__35630;
    wire N__35629;
    wire N__35628;
    wire N__35625;
    wire N__35616;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35604;
    wire N__35601;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35571;
    wire N__35570;
    wire N__35569;
    wire N__35568;
    wire N__35565;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35508;
    wire N__35505;
    wire N__35502;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35490;
    wire N__35487;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35475;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35463;
    wire N__35460;
    wire N__35457;
    wire N__35454;
    wire N__35451;
    wire N__35450;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35412;
    wire N__35409;
    wire N__35408;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35400;
    wire N__35397;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35384;
    wire N__35383;
    wire N__35380;
    wire N__35377;
    wire N__35374;
    wire N__35369;
    wire N__35366;
    wire N__35355;
    wire N__35354;
    wire N__35353;
    wire N__35352;
    wire N__35347;
    wire N__35342;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35321;
    wire N__35316;
    wire N__35313;
    wire N__35310;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35298;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35286;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35265;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35253;
    wire N__35250;
    wire N__35247;
    wire N__35244;
    wire N__35241;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35229;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35193;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35164;
    wire N__35163;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35142;
    wire N__35139;
    wire N__35138;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35118;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35058;
    wire N__35055;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35043;
    wire N__35040;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35016;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34986;
    wire N__34985;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34970;
    wire N__34965;
    wire N__34964;
    wire N__34959;
    wire N__34958;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34919;
    wire N__34918;
    wire N__34917;
    wire N__34916;
    wire N__34913;
    wire N__34904;
    wire N__34899;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34891;
    wire N__34890;
    wire N__34889;
    wire N__34884;
    wire N__34881;
    wire N__34876;
    wire N__34869;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34791;
    wire N__34790;
    wire N__34787;
    wire N__34784;
    wire N__34779;
    wire N__34776;
    wire N__34775;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34656;
    wire N__34653;
    wire N__34650;
    wire N__34647;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34626;
    wire N__34623;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34574;
    wire N__34573;
    wire N__34572;
    wire N__34571;
    wire N__34570;
    wire N__34569;
    wire N__34568;
    wire N__34567;
    wire N__34564;
    wire N__34563;
    wire N__34562;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34557;
    wire N__34556;
    wire N__34555;
    wire N__34554;
    wire N__34553;
    wire N__34552;
    wire N__34551;
    wire N__34548;
    wire N__34541;
    wire N__34532;
    wire N__34531;
    wire N__34530;
    wire N__34529;
    wire N__34528;
    wire N__34525;
    wire N__34516;
    wire N__34515;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34511;
    wire N__34510;
    wire N__34509;
    wire N__34508;
    wire N__34507;
    wire N__34506;
    wire N__34503;
    wire N__34502;
    wire N__34499;
    wire N__34492;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34474;
    wire N__34465;
    wire N__34460;
    wire N__34451;
    wire N__34442;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34396;
    wire N__34391;
    wire N__34386;
    wire N__34383;
    wire N__34378;
    wire N__34375;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34361;
    wire N__34358;
    wire N__34357;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34341;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34311;
    wire N__34310;
    wire N__34309;
    wire N__34308;
    wire N__34303;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34278;
    wire N__34275;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34265;
    wire N__34262;
    wire N__34259;
    wire N__34254;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34232;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34217;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34176;
    wire N__34173;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34158;
    wire N__34155;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34145;
    wire N__34140;
    wire N__34137;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34122;
    wire N__34119;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34104;
    wire N__34101;
    wire N__34100;
    wire N__34097;
    wire N__34094;
    wire N__34091;
    wire N__34086;
    wire N__34083;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34068;
    wire N__34065;
    wire N__34064;
    wire N__34061;
    wire N__34056;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34041;
    wire N__34038;
    wire N__34037;
    wire N__34034;
    wire N__34029;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33998;
    wire N__33995;
    wire N__33992;
    wire N__33989;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33957;
    wire N__33954;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33939;
    wire N__33936;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33921;
    wire N__33918;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33903;
    wire N__33900;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33828;
    wire N__33825;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33800;
    wire N__33795;
    wire N__33792;
    wire N__33791;
    wire N__33788;
    wire N__33785;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33717;
    wire N__33714;
    wire N__33711;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33675;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33432;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33380;
    wire N__33379;
    wire N__33376;
    wire N__33371;
    wire N__33366;
    wire N__33363;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33351;
    wire N__33348;
    wire N__33347;
    wire N__33344;
    wire N__33341;
    wire N__33340;
    wire N__33335;
    wire N__33332;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33314;
    wire N__33311;
    wire N__33310;
    wire N__33309;
    wire N__33308;
    wire N__33307;
    wire N__33306;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33294;
    wire N__33293;
    wire N__33292;
    wire N__33291;
    wire N__33288;
    wire N__33283;
    wire N__33278;
    wire N__33275;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33257;
    wire N__33252;
    wire N__33243;
    wire N__33242;
    wire N__33241;
    wire N__33240;
    wire N__33239;
    wire N__33238;
    wire N__33237;
    wire N__33236;
    wire N__33235;
    wire N__33234;
    wire N__33231;
    wire N__33230;
    wire N__33229;
    wire N__33228;
    wire N__33227;
    wire N__33226;
    wire N__33225;
    wire N__33224;
    wire N__33223;
    wire N__33216;
    wire N__33213;
    wire N__33204;
    wire N__33203;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33191;
    wire N__33190;
    wire N__33189;
    wire N__33188;
    wire N__33187;
    wire N__33186;
    wire N__33185;
    wire N__33184;
    wire N__33183;
    wire N__33182;
    wire N__33181;
    wire N__33180;
    wire N__33167;
    wire N__33164;
    wire N__33159;
    wire N__33154;
    wire N__33151;
    wire N__33146;
    wire N__33135;
    wire N__33132;
    wire N__33127;
    wire N__33122;
    wire N__33121;
    wire N__33120;
    wire N__33119;
    wire N__33118;
    wire N__33117;
    wire N__33114;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33088;
    wire N__33085;
    wire N__33078;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33062;
    wire N__33057;
    wire N__33042;
    wire N__33041;
    wire N__33040;
    wire N__33037;
    wire N__33036;
    wire N__33035;
    wire N__33034;
    wire N__33031;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33019;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33007;
    wire N__33004;
    wire N__33003;
    wire N__33000;
    wire N__32999;
    wire N__32998;
    wire N__32997;
    wire N__32996;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32961;
    wire N__32958;
    wire N__32949;
    wire N__32934;
    wire N__32931;
    wire N__32930;
    wire N__32927;
    wire N__32924;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32900;
    wire N__32899;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32866;
    wire N__32865;
    wire N__32864;
    wire N__32863;
    wire N__32862;
    wire N__32861;
    wire N__32860;
    wire N__32859;
    wire N__32858;
    wire N__32857;
    wire N__32856;
    wire N__32855;
    wire N__32854;
    wire N__32853;
    wire N__32852;
    wire N__32851;
    wire N__32850;
    wire N__32849;
    wire N__32848;
    wire N__32847;
    wire N__32846;
    wire N__32845;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32812;
    wire N__32803;
    wire N__32794;
    wire N__32785;
    wire N__32778;
    wire N__32769;
    wire N__32766;
    wire N__32765;
    wire N__32764;
    wire N__32763;
    wire N__32762;
    wire N__32761;
    wire N__32760;
    wire N__32759;
    wire N__32758;
    wire N__32751;
    wire N__32746;
    wire N__32743;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32717;
    wire N__32708;
    wire N__32703;
    wire N__32696;
    wire N__32685;
    wire N__32682;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32670;
    wire N__32669;
    wire N__32666;
    wire N__32663;
    wire N__32658;
    wire N__32655;
    wire N__32654;
    wire N__32651;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32599;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32582;
    wire N__32577;
    wire N__32574;
    wire N__32573;
    wire N__32570;
    wire N__32567;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32557;
    wire N__32554;
    wire N__32549;
    wire N__32544;
    wire N__32541;
    wire N__32540;
    wire N__32539;
    wire N__32536;
    wire N__32531;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32507;
    wire N__32504;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32487;
    wire N__32486;
    wire N__32483;
    wire N__32480;
    wire N__32479;
    wire N__32474;
    wire N__32471;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32429;
    wire N__32426;
    wire N__32423;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32384;
    wire N__32383;
    wire N__32380;
    wire N__32377;
    wire N__32374;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32344;
    wire N__32341;
    wire N__32336;
    wire N__32331;
    wire N__32328;
    wire N__32327;
    wire N__32326;
    wire N__32323;
    wire N__32322;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32295;
    wire N__32292;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32270;
    wire N__32267;
    wire N__32266;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32241;
    wire N__32238;
    wire N__32233;
    wire N__32230;
    wire N__32227;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32185;
    wire N__32182;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32168;
    wire N__32167;
    wire N__32164;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32153;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32108;
    wire N__32105;
    wire N__32102;
    wire N__32099;
    wire N__32096;
    wire N__32093;
    wire N__32092;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32080;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31994;
    wire N__31991;
    wire N__31988;
    wire N__31987;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31961;
    wire N__31958;
    wire N__31955;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31941;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31907;
    wire N__31904;
    wire N__31901;
    wire N__31900;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31886;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31867;
    wire N__31860;
    wire N__31857;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31847;
    wire N__31844;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31836;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31821;
    wire N__31818;
    wire N__31813;
    wire N__31810;
    wire N__31807;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31761;
    wire N__31760;
    wire N__31757;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31742;
    wire N__31739;
    wire N__31736;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31718;
    wire N__31717;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31707;
    wire N__31706;
    wire N__31701;
    wire N__31698;
    wire N__31693;
    wire N__31686;
    wire N__31683;
    wire N__31682;
    wire N__31679;
    wire N__31676;
    wire N__31673;
    wire N__31670;
    wire N__31667;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31649;
    wire N__31648;
    wire N__31645;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31613;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31589;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31567;
    wire N__31562;
    wire N__31559;
    wire N__31558;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31542;
    wire N__31541;
    wire N__31538;
    wire N__31537;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31524;
    wire N__31521;
    wire N__31516;
    wire N__31513;
    wire N__31506;
    wire N__31505;
    wire N__31504;
    wire N__31503;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31495;
    wire N__31494;
    wire N__31493;
    wire N__31490;
    wire N__31489;
    wire N__31480;
    wire N__31479;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31456;
    wire N__31453;
    wire N__31448;
    wire N__31443;
    wire N__31442;
    wire N__31441;
    wire N__31440;
    wire N__31439;
    wire N__31438;
    wire N__31437;
    wire N__31434;
    wire N__31433;
    wire N__31432;
    wire N__31431;
    wire N__31430;
    wire N__31429;
    wire N__31426;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31410;
    wire N__31401;
    wire N__31400;
    wire N__31399;
    wire N__31398;
    wire N__31397;
    wire N__31396;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31382;
    wire N__31377;
    wire N__31376;
    wire N__31373;
    wire N__31372;
    wire N__31371;
    wire N__31370;
    wire N__31359;
    wire N__31350;
    wire N__31347;
    wire N__31346;
    wire N__31345;
    wire N__31344;
    wire N__31341;
    wire N__31334;
    wire N__31331;
    wire N__31326;
    wire N__31323;
    wire N__31318;
    wire N__31305;
    wire N__31304;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31291;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31279;
    wire N__31272;
    wire N__31269;
    wire N__31268;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31236;
    wire N__31235;
    wire N__31232;
    wire N__31231;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31213;
    wire N__31210;
    wire N__31203;
    wire N__31200;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31188;
    wire N__31185;
    wire N__31184;
    wire N__31181;
    wire N__31178;
    wire N__31173;
    wire N__31172;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31155;
    wire N__31152;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31124;
    wire N__31123;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31112;
    wire N__31111;
    wire N__31110;
    wire N__31109;
    wire N__31108;
    wire N__31107;
    wire N__31106;
    wire N__31105;
    wire N__31104;
    wire N__31103;
    wire N__31100;
    wire N__31099;
    wire N__31094;
    wire N__31093;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31085;
    wire N__31082;
    wire N__31081;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31073;
    wire N__31072;
    wire N__31069;
    wire N__31068;
    wire N__31067;
    wire N__31066;
    wire N__31063;
    wire N__31058;
    wire N__31057;
    wire N__31056;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31044;
    wire N__31043;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31028;
    wire N__31019;
    wire N__31010;
    wire N__30999;
    wire N__30996;
    wire N__30987;
    wire N__30982;
    wire N__30977;
    wire N__30954;
    wire N__30951;
    wire N__30950;
    wire N__30949;
    wire N__30946;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30924;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30899;
    wire N__30896;
    wire N__30893;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30870;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30810;
    wire N__30807;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30786;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30762;
    wire N__30759;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30747;
    wire N__30744;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30686;
    wire N__30685;
    wire N__30684;
    wire N__30681;
    wire N__30678;
    wire N__30677;
    wire N__30674;
    wire N__30673;
    wire N__30672;
    wire N__30671;
    wire N__30670;
    wire N__30669;
    wire N__30668;
    wire N__30667;
    wire N__30666;
    wire N__30665;
    wire N__30664;
    wire N__30663;
    wire N__30662;
    wire N__30661;
    wire N__30658;
    wire N__30657;
    wire N__30656;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30644;
    wire N__30641;
    wire N__30634;
    wire N__30627;
    wire N__30616;
    wire N__30607;
    wire N__30604;
    wire N__30597;
    wire N__30582;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30570;
    wire N__30567;
    wire N__30566;
    wire N__30563;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30548;
    wire N__30545;
    wire N__30540;
    wire N__30539;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30494;
    wire N__30493;
    wire N__30490;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30468;
    wire N__30467;
    wire N__30464;
    wire N__30461;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30443;
    wire N__30442;
    wire N__30437;
    wire N__30434;
    wire N__30433;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30415;
    wire N__30408;
    wire N__30407;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30392;
    wire N__30391;
    wire N__30390;
    wire N__30389;
    wire N__30386;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30366;
    wire N__30363;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30351;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30323;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30305;
    wire N__30300;
    wire N__30297;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30279;
    wire N__30278;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30254;
    wire N__30253;
    wire N__30252;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30238;
    wire N__30233;
    wire N__30232;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30195;
    wire N__30194;
    wire N__30191;
    wire N__30190;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30155;
    wire N__30154;
    wire N__30151;
    wire N__30150;
    wire N__30149;
    wire N__30144;
    wire N__30141;
    wire N__30136;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30122;
    wire N__30119;
    wire N__30118;
    wire N__30115;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30094;
    wire N__30087;
    wire N__30084;
    wire N__30083;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30066;
    wire N__30065;
    wire N__30064;
    wire N__30063;
    wire N__30062;
    wire N__30059;
    wire N__30058;
    wire N__30057;
    wire N__30052;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30022;
    wire N__30009;
    wire N__30006;
    wire N__30005;
    wire N__30002;
    wire N__30001;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29985;
    wire N__29982;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29961;
    wire N__29960;
    wire N__29957;
    wire N__29952;
    wire N__29951;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29928;
    wire N__29925;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29907;
    wire N__29904;
    wire N__29901;
    wire N__29898;
    wire N__29895;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29885;
    wire N__29884;
    wire N__29881;
    wire N__29876;
    wire N__29871;
    wire N__29868;
    wire N__29867;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29851;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29814;
    wire N__29813;
    wire N__29810;
    wire N__29807;
    wire N__29806;
    wire N__29805;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29789;
    wire N__29784;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29721;
    wire N__29720;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29703;
    wire N__29700;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29687;
    wire N__29684;
    wire N__29681;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29652;
    wire N__29651;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29598;
    wire N__29597;
    wire N__29594;
    wire N__29591;
    wire N__29588;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29516;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29501;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29450;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29429;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29397;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29389;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29363;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29348;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29222;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29176;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29097;
    wire N__29094;
    wire N__29091;
    wire N__29090;
    wire N__29087;
    wire N__29084;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29066;
    wire N__29065;
    wire N__29064;
    wire N__29061;
    wire N__29058;
    wire N__29053;
    wire N__29046;
    wire N__29045;
    wire N__29042;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29024;
    wire N__29021;
    wire N__29016;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29003;
    wire N__29000;
    wire N__28999;
    wire N__28998;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28962;
    wire N__28957;
    wire N__28950;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28937;
    wire N__28934;
    wire N__28933;
    wire N__28930;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28889;
    wire N__28884;
    wire N__28883;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28869;
    wire N__28866;
    wire N__28865;
    wire N__28860;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28845;
    wire N__28842;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28828;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28812;
    wire N__28811;
    wire N__28808;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28793;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28776;
    wire N__28775;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28761;
    wire N__28760;
    wire N__28757;
    wire N__28754;
    wire N__28751;
    wire N__28748;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28736;
    wire N__28735;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28674;
    wire N__28671;
    wire N__28670;
    wire N__28667;
    wire N__28664;
    wire N__28659;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28626;
    wire N__28623;
    wire N__28622;
    wire N__28621;
    wire N__28620;
    wire N__28619;
    wire N__28618;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28598;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28575;
    wire N__28572;
    wire N__28571;
    wire N__28568;
    wire N__28565;
    wire N__28562;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28537;
    wire N__28532;
    wire N__28529;
    wire N__28526;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28507;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28491;
    wire N__28488;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28480;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28464;
    wire N__28461;
    wire N__28460;
    wire N__28459;
    wire N__28454;
    wire N__28451;
    wire N__28448;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28429;
    wire N__28424;
    wire N__28421;
    wire N__28418;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28395;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28366;
    wire N__28361;
    wire N__28358;
    wire N__28355;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28336;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28320;
    wire N__28317;
    wire N__28316;
    wire N__28311;
    wire N__28310;
    wire N__28307;
    wire N__28304;
    wire N__28301;
    wire N__28296;
    wire N__28293;
    wire N__28292;
    wire N__28291;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28255;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28211;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28175;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28163;
    wire N__28158;
    wire N__28155;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28140;
    wire N__28137;
    wire N__28136;
    wire N__28131;
    wire N__28130;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28116;
    wire N__28113;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28101;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28086;
    wire N__28083;
    wire N__28082;
    wire N__28079;
    wire N__28078;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28042;
    wire N__28037;
    wire N__28034;
    wire N__28031;
    wire N__28026;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27990;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27978;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27951;
    wire N__27948;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27938;
    wire N__27937;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27921;
    wire N__27918;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27882;
    wire N__27879;
    wire N__27878;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27864;
    wire N__27861;
    wire N__27860;
    wire N__27857;
    wire N__27854;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27839;
    wire N__27836;
    wire N__27833;
    wire N__27828;
    wire N__27825;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27815;
    wire N__27810;
    wire N__27807;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27795;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27783;
    wire N__27780;
    wire N__27779;
    wire N__27778;
    wire N__27773;
    wire N__27770;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27758;
    wire N__27755;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27744;
    wire N__27743;
    wire N__27742;
    wire N__27735;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27722;
    wire N__27719;
    wire N__27714;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27630;
    wire N__27629;
    wire N__27628;
    wire N__27627;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27608;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27570;
    wire N__27569;
    wire N__27566;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27550;
    wire N__27547;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27524;
    wire N__27523;
    wire N__27522;
    wire N__27521;
    wire N__27520;
    wire N__27519;
    wire N__27518;
    wire N__27517;
    wire N__27516;
    wire N__27515;
    wire N__27514;
    wire N__27513;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27502;
    wire N__27501;
    wire N__27500;
    wire N__27499;
    wire N__27498;
    wire N__27497;
    wire N__27496;
    wire N__27481;
    wire N__27478;
    wire N__27477;
    wire N__27476;
    wire N__27475;
    wire N__27474;
    wire N__27473;
    wire N__27470;
    wire N__27459;
    wire N__27454;
    wire N__27443;
    wire N__27440;
    wire N__27439;
    wire N__27438;
    wire N__27437;
    wire N__27436;
    wire N__27435;
    wire N__27434;
    wire N__27431;
    wire N__27420;
    wire N__27413;
    wire N__27408;
    wire N__27405;
    wire N__27394;
    wire N__27391;
    wire N__27386;
    wire N__27383;
    wire N__27372;
    wire N__27371;
    wire N__27370;
    wire N__27369;
    wire N__27362;
    wire N__27361;
    wire N__27360;
    wire N__27359;
    wire N__27358;
    wire N__27357;
    wire N__27356;
    wire N__27355;
    wire N__27354;
    wire N__27353;
    wire N__27352;
    wire N__27351;
    wire N__27350;
    wire N__27349;
    wire N__27348;
    wire N__27347;
    wire N__27346;
    wire N__27345;
    wire N__27344;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27318;
    wire N__27317;
    wire N__27316;
    wire N__27315;
    wire N__27314;
    wire N__27313;
    wire N__27312;
    wire N__27311;
    wire N__27296;
    wire N__27285;
    wire N__27278;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27263;
    wire N__27260;
    wire N__27249;
    wire N__27244;
    wire N__27241;
    wire N__27238;
    wire N__27233;
    wire N__27226;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27197;
    wire N__27196;
    wire N__27195;
    wire N__27192;
    wire N__27191;
    wire N__27190;
    wire N__27189;
    wire N__27188;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27177;
    wire N__27176;
    wire N__27175;
    wire N__27174;
    wire N__27171;
    wire N__27170;
    wire N__27169;
    wire N__27168;
    wire N__27167;
    wire N__27166;
    wire N__27165;
    wire N__27164;
    wire N__27163;
    wire N__27162;
    wire N__27161;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27140;
    wire N__27139;
    wire N__27138;
    wire N__27137;
    wire N__27134;
    wire N__27133;
    wire N__27132;
    wire N__27129;
    wire N__27128;
    wire N__27127;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27100;
    wire N__27085;
    wire N__27082;
    wire N__27071;
    wire N__27066;
    wire N__27055;
    wire N__27050;
    wire N__27043;
    wire N__27040;
    wire N__27027;
    wire N__27026;
    wire N__27023;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27009;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26983;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26948;
    wire N__26943;
    wire N__26940;
    wire N__26939;
    wire N__26934;
    wire N__26931;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26923;
    wire N__26922;
    wire N__26921;
    wire N__26916;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26898;
    wire N__26897;
    wire N__26896;
    wire N__26893;
    wire N__26892;
    wire N__26891;
    wire N__26886;
    wire N__26883;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26846;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26832;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26817;
    wire N__26812;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26729;
    wire N__26728;
    wire N__26727;
    wire N__26722;
    wire N__26717;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26683;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26659;
    wire N__26654;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26554;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26535;
    wire N__26532;
    wire N__26527;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26510;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26481;
    wire N__26478;
    wire N__26473;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26424;
    wire N__26421;
    wire N__26420;
    wire N__26417;
    wire N__26416;
    wire N__26415;
    wire N__26412;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26380;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26350;
    wire N__26349;
    wire N__26344;
    wire N__26339;
    wire N__26338;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26322;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26300;
    wire N__26299;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26268;
    wire N__26265;
    wire N__26260;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26197;
    wire N__26192;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26169;
    wire N__26168;
    wire N__26167;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26154;
    wire N__26151;
    wire N__26146;
    wire N__26143;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26106;
    wire N__26105;
    wire N__26102;
    wire N__26099;
    wire N__26094;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26024;
    wire N__26021;
    wire N__26020;
    wire N__26017;
    wire N__26014;
    wire N__26013;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__25998;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25929;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25917;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25905;
    wire N__25902;
    wire N__25899;
    wire N__25896;
    wire N__25895;
    wire N__25894;
    wire N__25891;
    wire N__25886;
    wire N__25881;
    wire N__25880;
    wire N__25877;
    wire N__25876;
    wire N__25873;
    wire N__25868;
    wire N__25863;
    wire N__25860;
    wire N__25857;
    wire N__25854;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25842;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25823;
    wire N__25822;
    wire N__25819;
    wire N__25814;
    wire N__25809;
    wire N__25808;
    wire N__25805;
    wire N__25800;
    wire N__25797;
    wire N__25794;
    wire N__25791;
    wire N__25790;
    wire N__25789;
    wire N__25786;
    wire N__25781;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25755;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25725;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25713;
    wire N__25710;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25679;
    wire N__25676;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25664;
    wire N__25663;
    wire N__25660;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25635;
    wire N__25632;
    wire N__25631;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25484;
    wire N__25481;
    wire N__25478;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25451;
    wire N__25448;
    wire N__25445;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25202;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25106;
    wire N__25105;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25070;
    wire N__25065;
    wire N__25062;
    wire N__25061;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24696;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24560;
    wire N__24559;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24496;
    wire N__24495;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24474;
    wire N__24473;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24351;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24339;
    wire N__24336;
    wire N__24335;
    wire N__24334;
    wire N__24333;
    wire N__24332;
    wire N__24329;
    wire N__24324;
    wire N__24319;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24269;
    wire N__24268;
    wire N__24267;
    wire N__24266;
    wire N__24265;
    wire N__24264;
    wire N__24263;
    wire N__24262;
    wire N__24261;
    wire N__24260;
    wire N__24259;
    wire N__24258;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24254;
    wire N__24253;
    wire N__24252;
    wire N__24251;
    wire N__24250;
    wire N__24249;
    wire N__24248;
    wire N__24247;
    wire N__24246;
    wire N__24245;
    wire N__24244;
    wire N__24243;
    wire N__24242;
    wire N__24241;
    wire N__24232;
    wire N__24223;
    wire N__24218;
    wire N__24209;
    wire N__24200;
    wire N__24191;
    wire N__24182;
    wire N__24173;
    wire N__24162;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24146;
    wire N__24145;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24113;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24053;
    wire N__24052;
    wire N__24051;
    wire N__24046;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24030;
    wire N__24029;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23988;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23942;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23921;
    wire N__23918;
    wire N__23911;
    wire N__23908;
    wire N__23901;
    wire N__23898;
    wire N__23897;
    wire N__23896;
    wire N__23895;
    wire N__23894;
    wire N__23893;
    wire N__23892;
    wire N__23891;
    wire N__23890;
    wire N__23887;
    wire N__23886;
    wire N__23883;
    wire N__23882;
    wire N__23879;
    wire N__23878;
    wire N__23875;
    wire N__23874;
    wire N__23871;
    wire N__23870;
    wire N__23867;
    wire N__23866;
    wire N__23863;
    wire N__23862;
    wire N__23861;
    wire N__23844;
    wire N__23827;
    wire N__23824;
    wire N__23823;
    wire N__23818;
    wire N__23813;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23801;
    wire N__23798;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23787;
    wire N__23786;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23772;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23729;
    wire N__23726;
    wire N__23725;
    wire N__23722;
    wire N__23721;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23706;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23645;
    wire N__23644;
    wire N__23643;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23625;
    wire N__23622;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23610;
    wire N__23609;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23562;
    wire N__23559;
    wire N__23558;
    wire N__23555;
    wire N__23554;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23542;
    wire N__23539;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23484;
    wire N__23483;
    wire N__23478;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23466;
    wire N__23465;
    wire N__23464;
    wire N__23459;
    wire N__23456;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23403;
    wire N__23400;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23241;
    wire N__23240;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23204;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23187;
    wire N__23184;
    wire N__23183;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23169;
    wire N__23166;
    wire N__23165;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23130;
    wire N__23127;
    wire N__23126;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23111;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23096;
    wire N__23091;
    wire N__23090;
    wire N__23089;
    wire N__23088;
    wire N__23087;
    wire N__23086;
    wire N__23083;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23068;
    wire N__23067;
    wire N__23066;
    wire N__23055;
    wire N__23050;
    wire N__23047;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23022;
    wire N__23019;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22977;
    wire N__22974;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22962;
    wire N__22959;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22947;
    wire N__22944;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22919;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22890;
    wire N__22887;
    wire N__22886;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22857;
    wire N__22854;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22846;
    wire N__22841;
    wire N__22838;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22823;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22811;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22793;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22781;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22769;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22703;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22657;
    wire N__22656;
    wire N__22651;
    wire N__22646;
    wire N__22641;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22625;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22610;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22589;
    wire N__22586;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22557;
    wire N__22556;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22539;
    wire N__22536;
    wire N__22535;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22518;
    wire N__22515;
    wire N__22514;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22497;
    wire N__22494;
    wire N__22493;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22476;
    wire N__22473;
    wire N__22472;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22455;
    wire N__22452;
    wire N__22451;
    wire N__22450;
    wire N__22449;
    wire N__22448;
    wire N__22447;
    wire N__22446;
    wire N__22445;
    wire N__22444;
    wire N__22443;
    wire N__22434;
    wire N__22429;
    wire N__22420;
    wire N__22413;
    wire N__22410;
    wire N__22409;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22361;
    wire N__22358;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22298;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22281;
    wire N__22278;
    wire N__22277;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22260;
    wire N__22257;
    wire N__22256;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22239;
    wire N__22236;
    wire N__22235;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22202;
    wire N__22201;
    wire N__22200;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22186;
    wire N__22185;
    wire N__22184;
    wire N__22181;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22154;
    wire N__22151;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22125;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22019;
    wire N__22018;
    wire N__22013;
    wire N__22010;
    wire N__22009;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21997;
    wire N__21990;
    wire N__21989;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21969;
    wire N__21966;
    wire N__21961;
    wire N__21958;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21947;
    wire N__21944;
    wire N__21943;
    wire N__21940;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21928;
    wire N__21927;
    wire N__21926;
    wire N__21925;
    wire N__21924;
    wire N__21923;
    wire N__21922;
    wire N__21921;
    wire N__21920;
    wire N__21919;
    wire N__21918;
    wire N__21917;
    wire N__21916;
    wire N__21915;
    wire N__21914;
    wire N__21913;
    wire N__21912;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21897;
    wire N__21894;
    wire N__21893;
    wire N__21892;
    wire N__21891;
    wire N__21888;
    wire N__21871;
    wire N__21856;
    wire N__21855;
    wire N__21854;
    wire N__21853;
    wire N__21852;
    wire N__21851;
    wire N__21848;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21826;
    wire N__21819;
    wire N__21812;
    wire N__21805;
    wire N__21802;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21784;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21761;
    wire N__21760;
    wire N__21759;
    wire N__21758;
    wire N__21753;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21741;
    wire N__21740;
    wire N__21737;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21725;
    wire N__21724;
    wire N__21723;
    wire N__21720;
    wire N__21713;
    wire N__21706;
    wire N__21703;
    wire N__21698;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21686;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21653;
    wire N__21650;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21620;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21605;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21548;
    wire N__21545;
    wire N__21542;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21528;
    wire N__21527;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21328;
    wire N__21327;
    wire N__21324;
    wire N__21323;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21312;
    wire N__21309;
    wire N__21304;
    wire N__21297;
    wire N__21296;
    wire N__21295;
    wire N__21294;
    wire N__21293;
    wire N__21292;
    wire N__21289;
    wire N__21284;
    wire N__21281;
    wire N__21274;
    wire N__21269;
    wire N__21266;
    wire N__21255;
    wire N__21252;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20978;
    wire N__20977;
    wire N__20972;
    wire N__20969;
    wire N__20968;
    wire N__20967;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20953;
    wire N__20952;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20735;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20723;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20708;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20600;
    wire N__20597;
    wire N__20594;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20556;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20541;
    wire N__20538;
    wire N__20535;
    wire N__20532;
    wire N__20529;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20412;
    wire N__20409;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20369;
    wire N__20368;
    wire N__20363;
    wire N__20360;
    wire N__20355;
    wire N__20354;
    wire N__20353;
    wire N__20348;
    wire N__20345;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20333;
    wire N__20332;
    wire N__20329;
    wire N__20324;
    wire N__20321;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20306;
    wire N__20305;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20287;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20265;
    wire N__20262;
    wire N__20261;
    wire N__20258;
    wire N__20255;
    wire N__20254;
    wire N__20251;
    wire N__20248;
    wire N__20245;
    wire N__20240;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20219;
    wire N__20218;
    wire N__20213;
    wire N__20210;
    wire N__20205;
    wire N__20204;
    wire N__20201;
    wire N__20200;
    wire N__20197;
    wire N__20192;
    wire N__20189;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20174;
    wire N__20169;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20121;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20111;
    wire N__20106;
    wire N__20105;
    wire N__20102;
    wire N__20099;
    wire N__20094;
    wire N__20093;
    wire N__20092;
    wire N__20087;
    wire N__20084;
    wire N__20079;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20071;
    wire N__20068;
    wire N__20063;
    wire N__20060;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19907;
    wire N__19906;
    wire N__19905;
    wire N__19902;
    wire N__19901;
    wire N__19898;
    wire N__19897;
    wire N__19894;
    wire N__19893;
    wire N__19892;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19862;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.N_149 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_15 ;
    wire bfn_1_14_0_;
    wire \pwm_generator_inst.un2_threshold_acc_2_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_18 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_19 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_20 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_21 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_22 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_23 ;
    wire bfn_1_15_0_;
    wire \pwm_generator_inst.un2_threshold_acc_2_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_24 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_2_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_1_25 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ;
    wire bfn_1_16_0_;
    wire un7_start_stop_0_a2;
    wire N_38_i_i;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire pwm_duty_input_7;
    wire pwm_duty_input_8;
    wire pwm_duty_input_9;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire pwm_duty_input_6;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_27_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_153 ;
    wire pwm_duty_input_5;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire pwm_duty_input_4;
    wire pwm_duty_input_3;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \current_shift_inst.PI_CTRL.N_154 ;
    wire \current_shift_inst.PI_CTRL.N_155 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.N_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_7 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_6 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_4 ;
    wire bfn_2_14_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ;
    wire bfn_2_15_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ;
    wire bfn_2_16_0_;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_16 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_17 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_0 ;
    wire bfn_2_18_0_;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_2 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_3 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_4 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_6 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_7 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_7 ;
    wire bfn_2_19_0_;
    wire \pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ;
    wire \pwm_generator_inst.un19_threshold_acc_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_8 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_1 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_3 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_3_11_0_;
    wire \pwm_generator_inst.thresholdZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.thresholdZ0Z_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.thresholdZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.thresholdZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_3_12_0_;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto9_2_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9 ;
    wire \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_0 ;
    wire bfn_3_15_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_8 ;
    wire bfn_3_16_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ;
    wire \pwm_generator_inst.un3_threshold_acc ;
    wire \pwm_generator_inst.un19_threshold_acc_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ;
    wire bfn_3_17_0_;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_5 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_0 ;
    wire \pwm_generator_inst.thresholdZ0Z_0 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_5 ;
    wire \pwm_generator_inst.thresholdZ0Z_9 ;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_9 ;
    wire \pwm_generator_inst.thresholdZ0Z_8 ;
    wire \pwm_generator_inst.N_16 ;
    wire N_19_1;
    wire \pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.threshold_ACCZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_53 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire bfn_4_12_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire bfn_4_13_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_acc_1_axb_10 ;
    wire il_max_comp2_c;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_5_9_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_5_10_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_5_11_0_;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_5_12_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire il_max_comp2_D1;
    wire il_min_comp2_c;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire il_min_comp2_D1;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa ;
    wire il_max_comp2_D2;
    wire il_min_comp2_D2;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.N_393_i ;
    wire \phase_controller_inst2.start_timer_hc_RNO_0_0 ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire start_stop_c;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire s4_phy_c;
    wire il_max_comp1_c;
    wire il_max_comp1_D1;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_72 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire bfn_8_15_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_8_16_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_8_17_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_8_18_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.N_394_i ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire bfn_8_23_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_8_24_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_8_25_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_8_26_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire s3_phy_c;
    wire il_min_comp1_c;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire delay_hc_input_c_g;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire bfn_9_9_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire bfn_9_10_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire bfn_9_11_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire bfn_9_12_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_30 ;
    wire bfn_9_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_ ;
    wire elapsed_time_ns_1_RNIUE3CP1_0_6_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ;
    wire elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire elapsed_time_ns_1_RNILGKEE1_0_4_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_342_i_cascade_ ;
    wire elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17 ;
    wire elapsed_time_ns_1_RNIFFC6P1_0_16;
    wire \phase_controller_inst1.stoper_hc.N_267_iZ0Z_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_267_iZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_9_22_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_9_23_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire bfn_9_24_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_9 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.N_71 ;
    wire \pll_inst.red_c_i ;
    wire \current_shift_inst.PI_CTRL.integrator_i_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un1_enablelt3_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_30 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.N_74 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_ ;
    wire elapsed_time_ns_1_RNIJEKEE1_0_2_cascade_;
    wire \phase_controller_inst1.stoper_hc.N_284 ;
    wire elapsed_time_ns_1_RNIJEKEE1_0_2;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire elapsed_time_ns_1_RNI1I3CP1_0_9;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_326_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_308 ;
    wire elapsed_time_ns_1_RNILGKEE1_0_4;
    wire elapsed_time_ns_1_RNIAMU8E1_0_27;
    wire elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_;
    wire elapsed_time_ns_1_RNI6IU8E1_0_23;
    wire elapsed_time_ns_1_RNI6IU8E1_0_23_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1 ;
    wire elapsed_time_ns_1_RNI9LU8E1_0_26;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_ ;
    wire elapsed_time_ns_1_RNI5HU8E1_0_22;
    wire elapsed_time_ns_1_RNI7JU8E1_0_24;
    wire elapsed_time_ns_1_RNIBNU8E1_0_28;
    wire \delay_measurement_inst.delay_hc_timer.N_365_clk_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_367 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_ ;
    wire elapsed_time_ns_1_RNIDDC6P1_0_14;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14 ;
    wire elapsed_time_ns_1_RNIMHKEE1_0_5;
    wire elapsed_time_ns_1_RNI5IV8E1_0_31_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire bfn_10_19_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_10_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_10_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_10_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.N_393_i_g ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire elapsed_time_ns_1_RNIGGC6P1_0_17;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ;
    wire bfn_11_8_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_8 ;
    wire bfn_11_9_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ;
    wire bfn_11_10_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ;
    wire bfn_11_11_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_31 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0 ;
    wire il_min_comp1_D1;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ;
    wire elapsed_time_ns_1_RNIRB3CP1_0_3;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3_cascade_ ;
    wire elapsed_time_ns_1_RNIOJKEE1_0_7;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ;
    wire elapsed_time_ns_1_RNI7IT8E1_0_15;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ;
    wire elapsed_time_ns_1_RNIUE3CP1_0_6;
    wire \phase_controller_inst1.stoper_hc.N_328_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire elapsed_time_ns_1_RNICOU8E1_0_29;
    wire elapsed_time_ns_1_RNI4GU8E1_0_21;
    wire elapsed_time_ns_1_RNICOU8E1_0_29_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire elapsed_time_ns_1_RNI8KU8E1_0_25;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire elapsed_time_ns_1_RNI2DT8E1_0_10_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire elapsed_time_ns_1_RNI4HV8E1_0_30;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_342_i ;
    wire elapsed_time_ns_1_RNIP93CP1_0_1;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ;
    wire elapsed_time_ns_1_RNI3FU8E1_0_20;
    wire elapsed_time_ns_1_RNI2DT8E1_0_10;
    wire elapsed_time_ns_1_RNI3ET8E1_0_11;
    wire elapsed_time_ns_1_RNI4FT8E1_0_12;
    wire elapsed_time_ns_1_RNI5GT8E1_0_13;
    wire \phase_controller_inst1.stoper_hc.N_316 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ;
    wire elapsed_time_ns_1_RNIHHC6P1_0_18;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNIPKKEE1_0_8;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17 ;
    wire \delay_measurement_inst.delay_hc_timer.N_365_clk ;
    wire elapsed_time_ns_1_RNIIIC6P1_0_19;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire state_ns_i_a2_1;
    wire \phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire il_max_comp1_D2;
    wire \phase_controller_inst1.hc_time_passed ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \delay_measurement_inst.delay_tr_timer.N_395_i ;
    wire delay_tr_input_c_g;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_12_10_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire bfn_12_11_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ;
    wire \phase_controller_inst1.stoper_hc.N_328 ;
    wire elapsed_time_ns_1_RNI5IV8E1_0_31;
    wire \phase_controller_inst1.stoper_hc.N_326 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_12_14_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_12_15_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire bfn_12_16_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire bfn_12_17_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_12_18_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_12_19_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_12_20_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire il_min_comp1_D2;
    wire T12_c;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire T01_c;
    wire bfn_13_7_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_13_8_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_13_9_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_13_10_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.control_input_18 ;
    wire bfn_13_11_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_13_12_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.control_input_31 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_13_16_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_13_17_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire bfn_13_18_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df22 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df22 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df20 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_inst1.time_passed_RNI7NN7 ;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \current_shift_inst.timer_s1.N_166_i ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire s1_phy_c;
    wire T23_c;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire state_3;
    wire T45_c;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire bfn_14_5_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_14_6_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_14_7_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_14_8_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_167_i ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.N_1460_i ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire bfn_14_14_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_14_15_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_14_16_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_14_17_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire bfn_14_21_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire bfn_14_22_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_14_23_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire bfn_14_24_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire bfn_15_8_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire bfn_15_9_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_15_10_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_15_11_0_;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire bfn_15_12_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ;
    wire bfn_15_13_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_15_14_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_15_15_0_;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.N_242_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire elapsed_time_ns_1_RNIQENQL1_0_9_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_15_20_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_15_21_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire bfn_15_22_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_df20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df28 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_26 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire elapsed_time_ns_1_RNISAHF91_0_13_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire elapsed_time_ns_1_RNIVEIF91_0_25;
    wire elapsed_time_ns_1_RNI1HIF91_0_27;
    wire elapsed_time_ns_1_RNIVEIF91_0_25_cascade_;
    wire elapsed_time_ns_1_RNISBIF91_0_22;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15_cascade_ ;
    wire elapsed_time_ns_1_RNI2IIF91_0_28;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ;
    wire elapsed_time_ns_1_RNI0GIF91_0_26;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ;
    wire \delay_measurement_inst.delay_tr9_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_390 ;
    wire \delay_measurement_inst.delay_tr_timer.N_390_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_391_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ;
    wire elapsed_time_ns_1_RNI6565M1_0_14_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14 ;
    wire \delay_measurement_inst.delay_tr_timer.N_382 ;
    wire \delay_measurement_inst.delay_tr_timer.N_382_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_371 ;
    wire \delay_measurement_inst.delay_tr_timer.N_356 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ;
    wire \delay_measurement_inst.delay_tr_timer.N_351_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_378 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4 ;
    wire \delay_measurement_inst.delay_tr_timer.N_360 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5 ;
    wire \phase_controller_inst1.stoper_tr.N_242 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire bfn_17_7_0_;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_17_8_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire bfn_17_9_0_;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire bfn_17_10_0_;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire bfn_17_11_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire bfn_17_12_0_;
    wire \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_17_13_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_17_14_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire elapsed_time_ns_1_RNIP7HF91_0_10;
    wire elapsed_time_ns_1_RNIR9HF91_0_12;
    wire elapsed_time_ns_1_RNISAHF91_0_13;
    wire elapsed_time_ns_1_RNIP7HF91_0_10_cascade_;
    wire elapsed_time_ns_1_RNI6565M1_0_14;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_ ;
    wire elapsed_time_ns_1_RNIQENQL1_0_9;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ;
    wire elapsed_time_ns_1_RNIK8NQL1_0_3_cascade_;
    wire \delay_measurement_inst.N_363 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ;
    wire elapsed_time_ns_1_RNIBA65M1_0_19_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ;
    wire elapsed_time_ns_1_RNIQ9IF91_0_20;
    wire elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_;
    wire elapsed_time_ns_1_RNIRAIF91_0_21;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15 ;
    wire elapsed_time_ns_1_RNIQ8HF91_0_11;
    wire elapsed_time_ns_1_RNI3JIF91_0_29;
    wire elapsed_time_ns_1_RNITCIF91_0_23;
    wire elapsed_time_ns_1_RNITCIF91_0_23_cascade_;
    wire elapsed_time_ns_1_RNIUDIF91_0_24;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ;
    wire elapsed_time_ns_1_RNIA965M1_0_18;
    wire elapsed_time_ns_1_RNICG2591_0_4_cascade_;
    wire elapsed_time_ns_1_RNI9865M1_0_17;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_ ;
    wire elapsed_time_ns_1_RNIRBJF91_0_30;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4 ;
    wire \delay_measurement_inst.delay_tr_timer.N_344 ;
    wire \delay_measurement_inst.delay_tr_timer.N_344_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_347 ;
    wire \delay_measurement_inst.delay_tr_timer.N_347_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_373_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_351 ;
    wire \delay_measurement_inst.delay_tr_timer.N_353 ;
    wire \delay_measurement_inst.delay_tr_timer.N_348 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire bfn_17_19_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire bfn_17_20_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_17_21_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_17_22_0_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.N_166_i_g ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire elapsed_time_ns_1_RNIDH2591_0_5;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire elapsed_time_ns_1_RNI8765M1_0_16;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire elapsed_time_ns_1_RNIK8NQL1_0_3;
    wire elapsed_time_ns_1_RNIAE2591_0_2;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_ ;
    wire elapsed_time_ns_1_RNINBNQL1_0_6_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ;
    wire elapsed_time_ns_1_RNIUCHF91_0_15;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire elapsed_time_ns_1_RNINBNQL1_0_6;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire bfn_18_18_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_18_19_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_18_20_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_18_21_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_396_i ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire elapsed_time_ns_1_RNIGK2591_0_8;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ;
    wire elapsed_time_ns_1_RNII6NQL1_0_1_cascade_;
    wire elapsed_time_ns_1_RNIBA65M1_0_19;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ;
    wire \delay_measurement_inst.delay_tr9 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1 ;
    wire elapsed_time_ns_1_RNIFJ2591_0_7;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire elapsed_time_ns_1_RNICG2591_0_4;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.N_395_i_g ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ;
    wire elapsed_time_ns_1_RNISCJF91_0_31;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ;
    wire elapsed_time_ns_1_RNII6NQL1_0_1;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__32022),
            .RESETB(N__25983),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__38282),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__38275),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__21925,N__21918,N__21923,N__21917,N__21924,N__21916,N__21926,N__21913,N__21919,N__21912,N__21920,N__21914,N__21921,N__21915,N__21922}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__38281,N__38278,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__38276,N__38280,N__38277,N__38279}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,\pwm_generator_inst.un2_threshold_acc_2_1_16 ,\pwm_generator_inst.un2_threshold_acc_2_1_15 ,\pwm_generator_inst.un2_threshold_acc_2_14 ,\pwm_generator_inst.un2_threshold_acc_2_13 ,\pwm_generator_inst.un2_threshold_acc_2_12 ,\pwm_generator_inst.un2_threshold_acc_2_11 ,\pwm_generator_inst.un2_threshold_acc_2_10 ,\pwm_generator_inst.un2_threshold_acc_2_9 ,\pwm_generator_inst.un2_threshold_acc_2_8 ,\pwm_generator_inst.un2_threshold_acc_2_7 ,\pwm_generator_inst.un2_threshold_acc_2_6 ,\pwm_generator_inst.un2_threshold_acc_2_5 ,\pwm_generator_inst.un2_threshold_acc_2_4 ,\pwm_generator_inst.un2_threshold_acc_2_3 ,\pwm_generator_inst.un2_threshold_acc_2_2 ,\pwm_generator_inst.un2_threshold_acc_2_1 ,\pwm_generator_inst.un2_threshold_acc_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_acc_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__38250),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__38243),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .ADDSUBBOT(),
            .A({dangling_wire_74,N__21853,N__21891,N__21854,N__21892,N__21855,N__20353,N__20368,N__20079,N__20337,N__20261,N__20218,N__20204,N__20105,N__20121,N__20136}),
            .C({dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90}),
            .B({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__38249,N__38246,dangling_wire_98,dangling_wire_99,dangling_wire_100,N__38244,N__38248,N__38245,N__38247}),
            .OHOLDTOP(),
            .O({dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_acc_1_25 ,\pwm_generator_inst.un2_threshold_acc_1_24 ,\pwm_generator_inst.un2_threshold_acc_1_23 ,\pwm_generator_inst.un2_threshold_acc_1_22 ,\pwm_generator_inst.un2_threshold_acc_1_21 ,\pwm_generator_inst.un2_threshold_acc_1_20 ,\pwm_generator_inst.un2_threshold_acc_1_19 ,\pwm_generator_inst.un2_threshold_acc_1_18 ,\pwm_generator_inst.un2_threshold_acc_1_17 ,\pwm_generator_inst.un2_threshold_acc_1_16 ,\pwm_generator_inst.un2_threshold_acc_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold_acc ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__50614),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__50616),
            .DIN(N__50615),
            .DOUT(N__50614),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__50616),
            .PADOUT(N__50615),
            .PADIN(N__50614),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__50605),
            .DIN(N__50604),
            .DOUT(N__50603),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__50605),
            .PADOUT(N__50604),
            .PADIN(N__50603),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34278),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__50596),
            .DIN(N__50595),
            .DOUT(N__50594),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__50596),
            .PADOUT(N__50595),
            .PADIN(N__50594),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__50587),
            .DIN(N__50586),
            .DOUT(N__50585),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__50587),
            .PADOUT(N__50586),
            .PADIN(N__50585),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__50578),
            .DIN(N__50577),
            .DOUT(N__50576),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__50578),
            .PADOUT(N__50577),
            .PADIN(N__50576),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35700),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__50569),
            .DIN(N__50568),
            .DOUT(N__50567),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__50569),
            .PADOUT(N__50568),
            .PADIN(N__50567),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21009),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__50560),
            .DIN(N__50559),
            .DOUT(N__50558),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__50560),
            .PADOUT(N__50559),
            .PADIN(N__50558),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__50551),
            .DIN(N__50550),
            .DOUT(N__50549),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__50551),
            .PADOUT(N__50550),
            .PADIN(N__50549),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35508),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__50542),
            .DIN(N__50541),
            .DOUT(N__50540),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__50542),
            .PADOUT(N__50541),
            .PADIN(N__50540),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34335),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__50533),
            .DIN(N__50532),
            .DOUT(N__50531),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__50533),
            .PADOUT(N__50532),
            .PADIN(N__50531),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__50524),
            .DIN(N__50523),
            .DOUT(N__50522),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__50524),
            .PADOUT(N__50523),
            .PADIN(N__50522),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35727),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__50515),
            .DIN(N__50514),
            .DOUT(N__50513),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__50515),
            .PADOUT(N__50514),
            .PADIN(N__50513),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23532),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__50506),
            .DIN(N__50505),
            .DOUT(N__50504),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__50506),
            .PADOUT(N__50505),
            .PADIN(N__50504),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__50497),
            .DIN(N__50496),
            .DOUT(N__50495),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__50497),
            .PADOUT(N__50496),
            .PADIN(N__50495),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24522),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__50488),
            .DIN(N__50487),
            .DOUT(N__50486),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__50488),
            .PADOUT(N__50487),
            .PADIN(N__50486),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35592),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__50479),
            .DIN(N__50478),
            .DOUT(N__50477),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__50479),
            .PADOUT(N__50478),
            .PADIN(N__50477),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__50470),
            .DIN(N__50469),
            .DOUT(N__50468),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__50470),
            .PADOUT(N__50469),
            .PADIN(N__50468),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11944 (
            .O(N__50451),
            .I(N__50448));
    LocalMux I__11943 (
            .O(N__50448),
            .I(N__50444));
    InMux I__11942 (
            .O(N__50447),
            .I(N__50441));
    Odrv4 I__11941 (
            .O(N__50444),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ));
    LocalMux I__11940 (
            .O(N__50441),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ));
    InMux I__11939 (
            .O(N__50436),
            .I(N__50433));
    LocalMux I__11938 (
            .O(N__50433),
            .I(N__50430));
    Odrv12 I__11937 (
            .O(N__50430),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__11936 (
            .O(N__50427),
            .I(N__50424));
    InMux I__11935 (
            .O(N__50424),
            .I(N__50421));
    LocalMux I__11934 (
            .O(N__50421),
            .I(N__50417));
    InMux I__11933 (
            .O(N__50420),
            .I(N__50413));
    Span4Mux_h I__11932 (
            .O(N__50417),
            .I(N__50410));
    InMux I__11931 (
            .O(N__50416),
            .I(N__50407));
    LocalMux I__11930 (
            .O(N__50413),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    Odrv4 I__11929 (
            .O(N__50410),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    LocalMux I__11928 (
            .O(N__50407),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    CascadeMux I__11927 (
            .O(N__50400),
            .I(N__50396));
    CascadeMux I__11926 (
            .O(N__50399),
            .I(N__50387));
    InMux I__11925 (
            .O(N__50396),
            .I(N__50376));
    InMux I__11924 (
            .O(N__50395),
            .I(N__50376));
    InMux I__11923 (
            .O(N__50394),
            .I(N__50376));
    InMux I__11922 (
            .O(N__50393),
            .I(N__50371));
    InMux I__11921 (
            .O(N__50392),
            .I(N__50371));
    InMux I__11920 (
            .O(N__50391),
            .I(N__50368));
    InMux I__11919 (
            .O(N__50390),
            .I(N__50363));
    InMux I__11918 (
            .O(N__50387),
            .I(N__50363));
    InMux I__11917 (
            .O(N__50386),
            .I(N__50360));
    InMux I__11916 (
            .O(N__50385),
            .I(N__50356));
    InMux I__11915 (
            .O(N__50384),
            .I(N__50353));
    CascadeMux I__11914 (
            .O(N__50383),
            .I(N__50350));
    LocalMux I__11913 (
            .O(N__50376),
            .I(N__50345));
    LocalMux I__11912 (
            .O(N__50371),
            .I(N__50342));
    LocalMux I__11911 (
            .O(N__50368),
            .I(N__50337));
    LocalMux I__11910 (
            .O(N__50363),
            .I(N__50337));
    LocalMux I__11909 (
            .O(N__50360),
            .I(N__50334));
    InMux I__11908 (
            .O(N__50359),
            .I(N__50331));
    LocalMux I__11907 (
            .O(N__50356),
            .I(N__50326));
    LocalMux I__11906 (
            .O(N__50353),
            .I(N__50326));
    InMux I__11905 (
            .O(N__50350),
            .I(N__50319));
    InMux I__11904 (
            .O(N__50349),
            .I(N__50319));
    InMux I__11903 (
            .O(N__50348),
            .I(N__50319));
    Span4Mux_v I__11902 (
            .O(N__50345),
            .I(N__50316));
    Span4Mux_v I__11901 (
            .O(N__50342),
            .I(N__50309));
    Span4Mux_v I__11900 (
            .O(N__50337),
            .I(N__50309));
    Span4Mux_v I__11899 (
            .O(N__50334),
            .I(N__50309));
    LocalMux I__11898 (
            .O(N__50331),
            .I(N__50306));
    Odrv4 I__11897 (
            .O(N__50326),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__11896 (
            .O(N__50319),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    Odrv4 I__11895 (
            .O(N__50316),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    Odrv4 I__11894 (
            .O(N__50309),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    Odrv4 I__11893 (
            .O(N__50306),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    InMux I__11892 (
            .O(N__50295),
            .I(N__50292));
    LocalMux I__11891 (
            .O(N__50292),
            .I(N__50289));
    Odrv12 I__11890 (
            .O(N__50289),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    CEMux I__11889 (
            .O(N__50286),
            .I(N__50281));
    CEMux I__11888 (
            .O(N__50285),
            .I(N__50273));
    CEMux I__11887 (
            .O(N__50284),
            .I(N__50270));
    LocalMux I__11886 (
            .O(N__50281),
            .I(N__50267));
    CEMux I__11885 (
            .O(N__50280),
            .I(N__50264));
    InMux I__11884 (
            .O(N__50279),
            .I(N__50252));
    InMux I__11883 (
            .O(N__50278),
            .I(N__50252));
    InMux I__11882 (
            .O(N__50277),
            .I(N__50252));
    CEMux I__11881 (
            .O(N__50276),
            .I(N__50234));
    LocalMux I__11880 (
            .O(N__50273),
            .I(N__50231));
    LocalMux I__11879 (
            .O(N__50270),
            .I(N__50226));
    Span4Mux_v I__11878 (
            .O(N__50267),
            .I(N__50226));
    LocalMux I__11877 (
            .O(N__50264),
            .I(N__50223));
    InMux I__11876 (
            .O(N__50263),
            .I(N__50214));
    InMux I__11875 (
            .O(N__50262),
            .I(N__50214));
    InMux I__11874 (
            .O(N__50261),
            .I(N__50214));
    InMux I__11873 (
            .O(N__50260),
            .I(N__50214));
    CEMux I__11872 (
            .O(N__50259),
            .I(N__50211));
    LocalMux I__11871 (
            .O(N__50252),
            .I(N__50208));
    InMux I__11870 (
            .O(N__50251),
            .I(N__50201));
    InMux I__11869 (
            .O(N__50250),
            .I(N__50201));
    InMux I__11868 (
            .O(N__50249),
            .I(N__50201));
    InMux I__11867 (
            .O(N__50248),
            .I(N__50192));
    InMux I__11866 (
            .O(N__50247),
            .I(N__50192));
    InMux I__11865 (
            .O(N__50246),
            .I(N__50192));
    InMux I__11864 (
            .O(N__50245),
            .I(N__50192));
    InMux I__11863 (
            .O(N__50244),
            .I(N__50183));
    InMux I__11862 (
            .O(N__50243),
            .I(N__50183));
    InMux I__11861 (
            .O(N__50242),
            .I(N__50183));
    InMux I__11860 (
            .O(N__50241),
            .I(N__50183));
    InMux I__11859 (
            .O(N__50240),
            .I(N__50174));
    InMux I__11858 (
            .O(N__50239),
            .I(N__50174));
    InMux I__11857 (
            .O(N__50238),
            .I(N__50174));
    InMux I__11856 (
            .O(N__50237),
            .I(N__50174));
    LocalMux I__11855 (
            .O(N__50234),
            .I(N__50171));
    Span4Mux_v I__11854 (
            .O(N__50231),
            .I(N__50167));
    Span4Mux_h I__11853 (
            .O(N__50226),
            .I(N__50164));
    Span4Mux_v I__11852 (
            .O(N__50223),
            .I(N__50153));
    LocalMux I__11851 (
            .O(N__50214),
            .I(N__50150));
    LocalMux I__11850 (
            .O(N__50211),
            .I(N__50137));
    Span4Mux_v I__11849 (
            .O(N__50208),
            .I(N__50137));
    LocalMux I__11848 (
            .O(N__50201),
            .I(N__50137));
    LocalMux I__11847 (
            .O(N__50192),
            .I(N__50137));
    LocalMux I__11846 (
            .O(N__50183),
            .I(N__50137));
    LocalMux I__11845 (
            .O(N__50174),
            .I(N__50137));
    Span4Mux_v I__11844 (
            .O(N__50171),
            .I(N__50134));
    InMux I__11843 (
            .O(N__50170),
            .I(N__50131));
    Span4Mux_h I__11842 (
            .O(N__50167),
            .I(N__50126));
    Span4Mux_h I__11841 (
            .O(N__50164),
            .I(N__50126));
    InMux I__11840 (
            .O(N__50163),
            .I(N__50117));
    InMux I__11839 (
            .O(N__50162),
            .I(N__50117));
    InMux I__11838 (
            .O(N__50161),
            .I(N__50117));
    InMux I__11837 (
            .O(N__50160),
            .I(N__50117));
    InMux I__11836 (
            .O(N__50159),
            .I(N__50108));
    InMux I__11835 (
            .O(N__50158),
            .I(N__50108));
    InMux I__11834 (
            .O(N__50157),
            .I(N__50108));
    InMux I__11833 (
            .O(N__50156),
            .I(N__50108));
    Span4Mux_h I__11832 (
            .O(N__50153),
            .I(N__50101));
    Span4Mux_v I__11831 (
            .O(N__50150),
            .I(N__50101));
    Span4Mux_v I__11830 (
            .O(N__50137),
            .I(N__50101));
    Span4Mux_h I__11829 (
            .O(N__50134),
            .I(N__50098));
    LocalMux I__11828 (
            .O(N__50131),
            .I(N__50087));
    Sp12to4 I__11827 (
            .O(N__50126),
            .I(N__50087));
    LocalMux I__11826 (
            .O(N__50117),
            .I(N__50087));
    LocalMux I__11825 (
            .O(N__50108),
            .I(N__50087));
    Sp12to4 I__11824 (
            .O(N__50101),
            .I(N__50087));
    Odrv4 I__11823 (
            .O(N__50098),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv12 I__11822 (
            .O(N__50087),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__11821 (
            .O(N__50082),
            .I(N__50078));
    CascadeMux I__11820 (
            .O(N__50081),
            .I(N__50075));
    LocalMux I__11819 (
            .O(N__50078),
            .I(N__50071));
    InMux I__11818 (
            .O(N__50075),
            .I(N__50068));
    InMux I__11817 (
            .O(N__50074),
            .I(N__50065));
    Odrv4 I__11816 (
            .O(N__50071),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__11815 (
            .O(N__50068),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__11814 (
            .O(N__50065),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    CascadeMux I__11813 (
            .O(N__50058),
            .I(N__50055));
    InMux I__11812 (
            .O(N__50055),
            .I(N__50051));
    InMux I__11811 (
            .O(N__50054),
            .I(N__50048));
    LocalMux I__11810 (
            .O(N__50051),
            .I(N__50045));
    LocalMux I__11809 (
            .O(N__50048),
            .I(N__50042));
    Odrv4 I__11808 (
            .O(N__50045),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    Odrv12 I__11807 (
            .O(N__50042),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__11806 (
            .O(N__50037),
            .I(N__50033));
    CascadeMux I__11805 (
            .O(N__50036),
            .I(N__50030));
    LocalMux I__11804 (
            .O(N__50033),
            .I(N__50026));
    InMux I__11803 (
            .O(N__50030),
            .I(N__50023));
    InMux I__11802 (
            .O(N__50029),
            .I(N__50020));
    Odrv4 I__11801 (
            .O(N__50026),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__11800 (
            .O(N__50023),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__11799 (
            .O(N__50020),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__11798 (
            .O(N__50013),
            .I(N__50010));
    LocalMux I__11797 (
            .O(N__50010),
            .I(N__50005));
    InMux I__11796 (
            .O(N__50009),
            .I(N__50000));
    InMux I__11795 (
            .O(N__50008),
            .I(N__50000));
    Span4Mux_v I__11794 (
            .O(N__50005),
            .I(N__49997));
    LocalMux I__11793 (
            .O(N__50000),
            .I(N__49994));
    Odrv4 I__11792 (
            .O(N__49997),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    Odrv12 I__11791 (
            .O(N__49994),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    CEMux I__11790 (
            .O(N__49989),
            .I(N__49974));
    CEMux I__11789 (
            .O(N__49988),
            .I(N__49974));
    CEMux I__11788 (
            .O(N__49987),
            .I(N__49974));
    CEMux I__11787 (
            .O(N__49986),
            .I(N__49974));
    CEMux I__11786 (
            .O(N__49985),
            .I(N__49974));
    GlobalMux I__11785 (
            .O(N__49974),
            .I(N__49971));
    gio2CtrlBuf I__11784 (
            .O(N__49971),
            .I(\delay_measurement_inst.delay_tr_timer.N_395_i_g ));
    InMux I__11783 (
            .O(N__49968),
            .I(N__49964));
    CascadeMux I__11782 (
            .O(N__49967),
            .I(N__49958));
    LocalMux I__11781 (
            .O(N__49964),
            .I(N__49955));
    InMux I__11780 (
            .O(N__49963),
            .I(N__49952));
    InMux I__11779 (
            .O(N__49962),
            .I(N__49948));
    InMux I__11778 (
            .O(N__49961),
            .I(N__49943));
    InMux I__11777 (
            .O(N__49958),
            .I(N__49943));
    Span4Mux_h I__11776 (
            .O(N__49955),
            .I(N__49940));
    LocalMux I__11775 (
            .O(N__49952),
            .I(N__49937));
    InMux I__11774 (
            .O(N__49951),
            .I(N__49934));
    LocalMux I__11773 (
            .O(N__49948),
            .I(N__49931));
    LocalMux I__11772 (
            .O(N__49943),
            .I(N__49928));
    Span4Mux_v I__11771 (
            .O(N__49940),
            .I(N__49925));
    Span12Mux_v I__11770 (
            .O(N__49937),
            .I(N__49922));
    LocalMux I__11769 (
            .O(N__49934),
            .I(N__49919));
    Span4Mux_v I__11768 (
            .O(N__49931),
            .I(N__49912));
    Span4Mux_v I__11767 (
            .O(N__49928),
            .I(N__49912));
    Span4Mux_h I__11766 (
            .O(N__49925),
            .I(N__49912));
    Odrv12 I__11765 (
            .O(N__49922),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv12 I__11764 (
            .O(N__49919),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__11763 (
            .O(N__49912),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    CascadeMux I__11762 (
            .O(N__49905),
            .I(N__49901));
    InMux I__11761 (
            .O(N__49904),
            .I(N__49897));
    InMux I__11760 (
            .O(N__49901),
            .I(N__49894));
    InMux I__11759 (
            .O(N__49900),
            .I(N__49890));
    LocalMux I__11758 (
            .O(N__49897),
            .I(N__49883));
    LocalMux I__11757 (
            .O(N__49894),
            .I(N__49880));
    InMux I__11756 (
            .O(N__49893),
            .I(N__49877));
    LocalMux I__11755 (
            .O(N__49890),
            .I(N__49871));
    InMux I__11754 (
            .O(N__49889),
            .I(N__49866));
    InMux I__11753 (
            .O(N__49888),
            .I(N__49866));
    CascadeMux I__11752 (
            .O(N__49887),
            .I(N__49857));
    CascadeMux I__11751 (
            .O(N__49886),
            .I(N__49854));
    Span4Mux_v I__11750 (
            .O(N__49883),
            .I(N__49849));
    Span4Mux_v I__11749 (
            .O(N__49880),
            .I(N__49849));
    LocalMux I__11748 (
            .O(N__49877),
            .I(N__49846));
    CascadeMux I__11747 (
            .O(N__49876),
            .I(N__49842));
    CascadeMux I__11746 (
            .O(N__49875),
            .I(N__49836));
    InMux I__11745 (
            .O(N__49874),
            .I(N__49833));
    Span4Mux_h I__11744 (
            .O(N__49871),
            .I(N__49828));
    LocalMux I__11743 (
            .O(N__49866),
            .I(N__49828));
    CascadeMux I__11742 (
            .O(N__49865),
            .I(N__49825));
    CascadeMux I__11741 (
            .O(N__49864),
            .I(N__49822));
    InMux I__11740 (
            .O(N__49863),
            .I(N__49806));
    InMux I__11739 (
            .O(N__49862),
            .I(N__49806));
    InMux I__11738 (
            .O(N__49861),
            .I(N__49806));
    InMux I__11737 (
            .O(N__49860),
            .I(N__49801));
    InMux I__11736 (
            .O(N__49857),
            .I(N__49801));
    InMux I__11735 (
            .O(N__49854),
            .I(N__49798));
    Span4Mux_h I__11734 (
            .O(N__49849),
            .I(N__49795));
    Span4Mux_h I__11733 (
            .O(N__49846),
            .I(N__49792));
    InMux I__11732 (
            .O(N__49845),
            .I(N__49783));
    InMux I__11731 (
            .O(N__49842),
            .I(N__49783));
    InMux I__11730 (
            .O(N__49841),
            .I(N__49783));
    InMux I__11729 (
            .O(N__49840),
            .I(N__49783));
    InMux I__11728 (
            .O(N__49839),
            .I(N__49778));
    InMux I__11727 (
            .O(N__49836),
            .I(N__49778));
    LocalMux I__11726 (
            .O(N__49833),
            .I(N__49775));
    Span4Mux_v I__11725 (
            .O(N__49828),
            .I(N__49772));
    InMux I__11724 (
            .O(N__49825),
            .I(N__49761));
    InMux I__11723 (
            .O(N__49822),
            .I(N__49761));
    InMux I__11722 (
            .O(N__49821),
            .I(N__49761));
    InMux I__11721 (
            .O(N__49820),
            .I(N__49761));
    InMux I__11720 (
            .O(N__49819),
            .I(N__49761));
    InMux I__11719 (
            .O(N__49818),
            .I(N__49758));
    InMux I__11718 (
            .O(N__49817),
            .I(N__49755));
    InMux I__11717 (
            .O(N__49816),
            .I(N__49746));
    InMux I__11716 (
            .O(N__49815),
            .I(N__49746));
    InMux I__11715 (
            .O(N__49814),
            .I(N__49746));
    InMux I__11714 (
            .O(N__49813),
            .I(N__49746));
    LocalMux I__11713 (
            .O(N__49806),
            .I(N__49743));
    LocalMux I__11712 (
            .O(N__49801),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__11711 (
            .O(N__49798),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__11710 (
            .O(N__49795),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__11709 (
            .O(N__49792),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__11708 (
            .O(N__49783),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__11707 (
            .O(N__49778),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__11706 (
            .O(N__49775),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__11705 (
            .O(N__49772),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__11704 (
            .O(N__49761),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__11703 (
            .O(N__49758),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__11702 (
            .O(N__49755),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__11701 (
            .O(N__49746),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__11700 (
            .O(N__49743),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    InMux I__11699 (
            .O(N__49716),
            .I(N__49712));
    InMux I__11698 (
            .O(N__49715),
            .I(N__49706));
    LocalMux I__11697 (
            .O(N__49712),
            .I(N__49702));
    CascadeMux I__11696 (
            .O(N__49711),
            .I(N__49697));
    CascadeMux I__11695 (
            .O(N__49710),
            .I(N__49693));
    CascadeMux I__11694 (
            .O(N__49709),
            .I(N__49687));
    LocalMux I__11693 (
            .O(N__49706),
            .I(N__49675));
    InMux I__11692 (
            .O(N__49705),
            .I(N__49672));
    Span4Mux_h I__11691 (
            .O(N__49702),
            .I(N__49669));
    InMux I__11690 (
            .O(N__49701),
            .I(N__49666));
    InMux I__11689 (
            .O(N__49700),
            .I(N__49663));
    InMux I__11688 (
            .O(N__49697),
            .I(N__49650));
    InMux I__11687 (
            .O(N__49696),
            .I(N__49650));
    InMux I__11686 (
            .O(N__49693),
            .I(N__49650));
    InMux I__11685 (
            .O(N__49692),
            .I(N__49650));
    InMux I__11684 (
            .O(N__49691),
            .I(N__49650));
    InMux I__11683 (
            .O(N__49690),
            .I(N__49650));
    InMux I__11682 (
            .O(N__49687),
            .I(N__49645));
    InMux I__11681 (
            .O(N__49686),
            .I(N__49645));
    InMux I__11680 (
            .O(N__49685),
            .I(N__49634));
    InMux I__11679 (
            .O(N__49684),
            .I(N__49634));
    InMux I__11678 (
            .O(N__49683),
            .I(N__49634));
    InMux I__11677 (
            .O(N__49682),
            .I(N__49634));
    InMux I__11676 (
            .O(N__49681),
            .I(N__49634));
    InMux I__11675 (
            .O(N__49680),
            .I(N__49627));
    InMux I__11674 (
            .O(N__49679),
            .I(N__49627));
    InMux I__11673 (
            .O(N__49678),
            .I(N__49627));
    Odrv12 I__11672 (
            .O(N__49675),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__11671 (
            .O(N__49672),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    Odrv4 I__11670 (
            .O(N__49669),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__11669 (
            .O(N__49666),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__11668 (
            .O(N__49663),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__11667 (
            .O(N__49650),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__11666 (
            .O(N__49645),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__11665 (
            .O(N__49634),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__11664 (
            .O(N__49627),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    CascadeMux I__11663 (
            .O(N__49608),
            .I(N__49603));
    CascadeMux I__11662 (
            .O(N__49607),
            .I(N__49600));
    InMux I__11661 (
            .O(N__49606),
            .I(N__49589));
    InMux I__11660 (
            .O(N__49603),
            .I(N__49589));
    InMux I__11659 (
            .O(N__49600),
            .I(N__49589));
    CascadeMux I__11658 (
            .O(N__49599),
            .I(N__49586));
    CascadeMux I__11657 (
            .O(N__49598),
            .I(N__49571));
    CascadeMux I__11656 (
            .O(N__49597),
            .I(N__49568));
    InMux I__11655 (
            .O(N__49596),
            .I(N__49561));
    LocalMux I__11654 (
            .O(N__49589),
            .I(N__49558));
    InMux I__11653 (
            .O(N__49586),
            .I(N__49545));
    InMux I__11652 (
            .O(N__49585),
            .I(N__49545));
    InMux I__11651 (
            .O(N__49584),
            .I(N__49545));
    InMux I__11650 (
            .O(N__49583),
            .I(N__49545));
    InMux I__11649 (
            .O(N__49582),
            .I(N__49545));
    InMux I__11648 (
            .O(N__49581),
            .I(N__49545));
    InMux I__11647 (
            .O(N__49580),
            .I(N__49542));
    CascadeMux I__11646 (
            .O(N__49579),
            .I(N__49539));
    InMux I__11645 (
            .O(N__49578),
            .I(N__49534));
    InMux I__11644 (
            .O(N__49577),
            .I(N__49527));
    InMux I__11643 (
            .O(N__49576),
            .I(N__49527));
    InMux I__11642 (
            .O(N__49575),
            .I(N__49527));
    InMux I__11641 (
            .O(N__49574),
            .I(N__49524));
    InMux I__11640 (
            .O(N__49571),
            .I(N__49517));
    InMux I__11639 (
            .O(N__49568),
            .I(N__49517));
    InMux I__11638 (
            .O(N__49567),
            .I(N__49517));
    InMux I__11637 (
            .O(N__49566),
            .I(N__49510));
    InMux I__11636 (
            .O(N__49565),
            .I(N__49510));
    InMux I__11635 (
            .O(N__49564),
            .I(N__49510));
    LocalMux I__11634 (
            .O(N__49561),
            .I(N__49507));
    Span4Mux_v I__11633 (
            .O(N__49558),
            .I(N__49502));
    LocalMux I__11632 (
            .O(N__49545),
            .I(N__49502));
    LocalMux I__11631 (
            .O(N__49542),
            .I(N__49499));
    InMux I__11630 (
            .O(N__49539),
            .I(N__49491));
    InMux I__11629 (
            .O(N__49538),
            .I(N__49491));
    InMux I__11628 (
            .O(N__49537),
            .I(N__49491));
    LocalMux I__11627 (
            .O(N__49534),
            .I(N__49486));
    LocalMux I__11626 (
            .O(N__49527),
            .I(N__49486));
    LocalMux I__11625 (
            .O(N__49524),
            .I(N__49483));
    LocalMux I__11624 (
            .O(N__49517),
            .I(N__49480));
    LocalMux I__11623 (
            .O(N__49510),
            .I(N__49475));
    Span4Mux_v I__11622 (
            .O(N__49507),
            .I(N__49475));
    Span4Mux_h I__11621 (
            .O(N__49502),
            .I(N__49470));
    Span4Mux_h I__11620 (
            .O(N__49499),
            .I(N__49470));
    CascadeMux I__11619 (
            .O(N__49498),
            .I(N__49461));
    LocalMux I__11618 (
            .O(N__49491),
            .I(N__49455));
    Span4Mux_v I__11617 (
            .O(N__49486),
            .I(N__49452));
    Span4Mux_v I__11616 (
            .O(N__49483),
            .I(N__49446));
    Span4Mux_v I__11615 (
            .O(N__49480),
            .I(N__49446));
    Sp12to4 I__11614 (
            .O(N__49475),
            .I(N__49441));
    Sp12to4 I__11613 (
            .O(N__49470),
            .I(N__49441));
    InMux I__11612 (
            .O(N__49469),
            .I(N__49432));
    InMux I__11611 (
            .O(N__49468),
            .I(N__49432));
    InMux I__11610 (
            .O(N__49467),
            .I(N__49432));
    InMux I__11609 (
            .O(N__49466),
            .I(N__49432));
    InMux I__11608 (
            .O(N__49465),
            .I(N__49427));
    InMux I__11607 (
            .O(N__49464),
            .I(N__49427));
    InMux I__11606 (
            .O(N__49461),
            .I(N__49424));
    InMux I__11605 (
            .O(N__49460),
            .I(N__49421));
    InMux I__11604 (
            .O(N__49459),
            .I(N__49416));
    InMux I__11603 (
            .O(N__49458),
            .I(N__49416));
    Span4Mux_h I__11602 (
            .O(N__49455),
            .I(N__49411));
    Span4Mux_h I__11601 (
            .O(N__49452),
            .I(N__49411));
    InMux I__11600 (
            .O(N__49451),
            .I(N__49408));
    Sp12to4 I__11599 (
            .O(N__49446),
            .I(N__49401));
    Span12Mux_v I__11598 (
            .O(N__49441),
            .I(N__49401));
    LocalMux I__11597 (
            .O(N__49432),
            .I(N__49401));
    LocalMux I__11596 (
            .O(N__49427),
            .I(N__49398));
    LocalMux I__11595 (
            .O(N__49424),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__11594 (
            .O(N__49421),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__11593 (
            .O(N__49416),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__11592 (
            .O(N__49411),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__11591 (
            .O(N__49408),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv12 I__11590 (
            .O(N__49401),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__11589 (
            .O(N__49398),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    InMux I__11588 (
            .O(N__49383),
            .I(N__49378));
    InMux I__11587 (
            .O(N__49382),
            .I(N__49375));
    InMux I__11586 (
            .O(N__49381),
            .I(N__49369));
    LocalMux I__11585 (
            .O(N__49378),
            .I(N__49361));
    LocalMux I__11584 (
            .O(N__49375),
            .I(N__49358));
    InMux I__11583 (
            .O(N__49374),
            .I(N__49351));
    InMux I__11582 (
            .O(N__49373),
            .I(N__49351));
    InMux I__11581 (
            .O(N__49372),
            .I(N__49351));
    LocalMux I__11580 (
            .O(N__49369),
            .I(N__49348));
    InMux I__11579 (
            .O(N__49368),
            .I(N__49343));
    InMux I__11578 (
            .O(N__49367),
            .I(N__49343));
    InMux I__11577 (
            .O(N__49366),
            .I(N__49336));
    InMux I__11576 (
            .O(N__49365),
            .I(N__49336));
    InMux I__11575 (
            .O(N__49364),
            .I(N__49336));
    Span4Mux_v I__11574 (
            .O(N__49361),
            .I(N__49331));
    Span4Mux_h I__11573 (
            .O(N__49358),
            .I(N__49331));
    LocalMux I__11572 (
            .O(N__49351),
            .I(N__49326));
    Span4Mux_h I__11571 (
            .O(N__49348),
            .I(N__49326));
    LocalMux I__11570 (
            .O(N__49343),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__11569 (
            .O(N__49336),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    Odrv4 I__11568 (
            .O(N__49331),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    Odrv4 I__11567 (
            .O(N__49326),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    InMux I__11566 (
            .O(N__49317),
            .I(N__49312));
    InMux I__11565 (
            .O(N__49316),
            .I(N__49309));
    InMux I__11564 (
            .O(N__49315),
            .I(N__49306));
    LocalMux I__11563 (
            .O(N__49312),
            .I(elapsed_time_ns_1_RNII6NQL1_0_1));
    LocalMux I__11562 (
            .O(N__49309),
            .I(elapsed_time_ns_1_RNII6NQL1_0_1));
    LocalMux I__11561 (
            .O(N__49306),
            .I(elapsed_time_ns_1_RNII6NQL1_0_1));
    CascadeMux I__11560 (
            .O(N__49299),
            .I(N__49295));
    InMux I__11559 (
            .O(N__49298),
            .I(N__49292));
    InMux I__11558 (
            .O(N__49295),
            .I(N__49289));
    LocalMux I__11557 (
            .O(N__49292),
            .I(N__49284));
    LocalMux I__11556 (
            .O(N__49289),
            .I(N__49284));
    Odrv4 I__11555 (
            .O(N__49284),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ));
    CascadeMux I__11554 (
            .O(N__49281),
            .I(N__49277));
    InMux I__11553 (
            .O(N__49280),
            .I(N__49274));
    InMux I__11552 (
            .O(N__49277),
            .I(N__49271));
    LocalMux I__11551 (
            .O(N__49274),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ));
    LocalMux I__11550 (
            .O(N__49271),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ));
    InMux I__11549 (
            .O(N__49266),
            .I(N__49263));
    LocalMux I__11548 (
            .O(N__49263),
            .I(N__49260));
    Span4Mux_h I__11547 (
            .O(N__49260),
            .I(N__49257));
    Span4Mux_v I__11546 (
            .O(N__49257),
            .I(N__49254));
    Odrv4 I__11545 (
            .O(N__49254),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    ClkMux I__11544 (
            .O(N__49251),
            .I(N__48825));
    ClkMux I__11543 (
            .O(N__49250),
            .I(N__48825));
    ClkMux I__11542 (
            .O(N__49249),
            .I(N__48825));
    ClkMux I__11541 (
            .O(N__49248),
            .I(N__48825));
    ClkMux I__11540 (
            .O(N__49247),
            .I(N__48825));
    ClkMux I__11539 (
            .O(N__49246),
            .I(N__48825));
    ClkMux I__11538 (
            .O(N__49245),
            .I(N__48825));
    ClkMux I__11537 (
            .O(N__49244),
            .I(N__48825));
    ClkMux I__11536 (
            .O(N__49243),
            .I(N__48825));
    ClkMux I__11535 (
            .O(N__49242),
            .I(N__48825));
    ClkMux I__11534 (
            .O(N__49241),
            .I(N__48825));
    ClkMux I__11533 (
            .O(N__49240),
            .I(N__48825));
    ClkMux I__11532 (
            .O(N__49239),
            .I(N__48825));
    ClkMux I__11531 (
            .O(N__49238),
            .I(N__48825));
    ClkMux I__11530 (
            .O(N__49237),
            .I(N__48825));
    ClkMux I__11529 (
            .O(N__49236),
            .I(N__48825));
    ClkMux I__11528 (
            .O(N__49235),
            .I(N__48825));
    ClkMux I__11527 (
            .O(N__49234),
            .I(N__48825));
    ClkMux I__11526 (
            .O(N__49233),
            .I(N__48825));
    ClkMux I__11525 (
            .O(N__49232),
            .I(N__48825));
    ClkMux I__11524 (
            .O(N__49231),
            .I(N__48825));
    ClkMux I__11523 (
            .O(N__49230),
            .I(N__48825));
    ClkMux I__11522 (
            .O(N__49229),
            .I(N__48825));
    ClkMux I__11521 (
            .O(N__49228),
            .I(N__48825));
    ClkMux I__11520 (
            .O(N__49227),
            .I(N__48825));
    ClkMux I__11519 (
            .O(N__49226),
            .I(N__48825));
    ClkMux I__11518 (
            .O(N__49225),
            .I(N__48825));
    ClkMux I__11517 (
            .O(N__49224),
            .I(N__48825));
    ClkMux I__11516 (
            .O(N__49223),
            .I(N__48825));
    ClkMux I__11515 (
            .O(N__49222),
            .I(N__48825));
    ClkMux I__11514 (
            .O(N__49221),
            .I(N__48825));
    ClkMux I__11513 (
            .O(N__49220),
            .I(N__48825));
    ClkMux I__11512 (
            .O(N__49219),
            .I(N__48825));
    ClkMux I__11511 (
            .O(N__49218),
            .I(N__48825));
    ClkMux I__11510 (
            .O(N__49217),
            .I(N__48825));
    ClkMux I__11509 (
            .O(N__49216),
            .I(N__48825));
    ClkMux I__11508 (
            .O(N__49215),
            .I(N__48825));
    ClkMux I__11507 (
            .O(N__49214),
            .I(N__48825));
    ClkMux I__11506 (
            .O(N__49213),
            .I(N__48825));
    ClkMux I__11505 (
            .O(N__49212),
            .I(N__48825));
    ClkMux I__11504 (
            .O(N__49211),
            .I(N__48825));
    ClkMux I__11503 (
            .O(N__49210),
            .I(N__48825));
    ClkMux I__11502 (
            .O(N__49209),
            .I(N__48825));
    ClkMux I__11501 (
            .O(N__49208),
            .I(N__48825));
    ClkMux I__11500 (
            .O(N__49207),
            .I(N__48825));
    ClkMux I__11499 (
            .O(N__49206),
            .I(N__48825));
    ClkMux I__11498 (
            .O(N__49205),
            .I(N__48825));
    ClkMux I__11497 (
            .O(N__49204),
            .I(N__48825));
    ClkMux I__11496 (
            .O(N__49203),
            .I(N__48825));
    ClkMux I__11495 (
            .O(N__49202),
            .I(N__48825));
    ClkMux I__11494 (
            .O(N__49201),
            .I(N__48825));
    ClkMux I__11493 (
            .O(N__49200),
            .I(N__48825));
    ClkMux I__11492 (
            .O(N__49199),
            .I(N__48825));
    ClkMux I__11491 (
            .O(N__49198),
            .I(N__48825));
    ClkMux I__11490 (
            .O(N__49197),
            .I(N__48825));
    ClkMux I__11489 (
            .O(N__49196),
            .I(N__48825));
    ClkMux I__11488 (
            .O(N__49195),
            .I(N__48825));
    ClkMux I__11487 (
            .O(N__49194),
            .I(N__48825));
    ClkMux I__11486 (
            .O(N__49193),
            .I(N__48825));
    ClkMux I__11485 (
            .O(N__49192),
            .I(N__48825));
    ClkMux I__11484 (
            .O(N__49191),
            .I(N__48825));
    ClkMux I__11483 (
            .O(N__49190),
            .I(N__48825));
    ClkMux I__11482 (
            .O(N__49189),
            .I(N__48825));
    ClkMux I__11481 (
            .O(N__49188),
            .I(N__48825));
    ClkMux I__11480 (
            .O(N__49187),
            .I(N__48825));
    ClkMux I__11479 (
            .O(N__49186),
            .I(N__48825));
    ClkMux I__11478 (
            .O(N__49185),
            .I(N__48825));
    ClkMux I__11477 (
            .O(N__49184),
            .I(N__48825));
    ClkMux I__11476 (
            .O(N__49183),
            .I(N__48825));
    ClkMux I__11475 (
            .O(N__49182),
            .I(N__48825));
    ClkMux I__11474 (
            .O(N__49181),
            .I(N__48825));
    ClkMux I__11473 (
            .O(N__49180),
            .I(N__48825));
    ClkMux I__11472 (
            .O(N__49179),
            .I(N__48825));
    ClkMux I__11471 (
            .O(N__49178),
            .I(N__48825));
    ClkMux I__11470 (
            .O(N__49177),
            .I(N__48825));
    ClkMux I__11469 (
            .O(N__49176),
            .I(N__48825));
    ClkMux I__11468 (
            .O(N__49175),
            .I(N__48825));
    ClkMux I__11467 (
            .O(N__49174),
            .I(N__48825));
    ClkMux I__11466 (
            .O(N__49173),
            .I(N__48825));
    ClkMux I__11465 (
            .O(N__49172),
            .I(N__48825));
    ClkMux I__11464 (
            .O(N__49171),
            .I(N__48825));
    ClkMux I__11463 (
            .O(N__49170),
            .I(N__48825));
    ClkMux I__11462 (
            .O(N__49169),
            .I(N__48825));
    ClkMux I__11461 (
            .O(N__49168),
            .I(N__48825));
    ClkMux I__11460 (
            .O(N__49167),
            .I(N__48825));
    ClkMux I__11459 (
            .O(N__49166),
            .I(N__48825));
    ClkMux I__11458 (
            .O(N__49165),
            .I(N__48825));
    ClkMux I__11457 (
            .O(N__49164),
            .I(N__48825));
    ClkMux I__11456 (
            .O(N__49163),
            .I(N__48825));
    ClkMux I__11455 (
            .O(N__49162),
            .I(N__48825));
    ClkMux I__11454 (
            .O(N__49161),
            .I(N__48825));
    ClkMux I__11453 (
            .O(N__49160),
            .I(N__48825));
    ClkMux I__11452 (
            .O(N__49159),
            .I(N__48825));
    ClkMux I__11451 (
            .O(N__49158),
            .I(N__48825));
    ClkMux I__11450 (
            .O(N__49157),
            .I(N__48825));
    ClkMux I__11449 (
            .O(N__49156),
            .I(N__48825));
    ClkMux I__11448 (
            .O(N__49155),
            .I(N__48825));
    ClkMux I__11447 (
            .O(N__49154),
            .I(N__48825));
    ClkMux I__11446 (
            .O(N__49153),
            .I(N__48825));
    ClkMux I__11445 (
            .O(N__49152),
            .I(N__48825));
    ClkMux I__11444 (
            .O(N__49151),
            .I(N__48825));
    ClkMux I__11443 (
            .O(N__49150),
            .I(N__48825));
    ClkMux I__11442 (
            .O(N__49149),
            .I(N__48825));
    ClkMux I__11441 (
            .O(N__49148),
            .I(N__48825));
    ClkMux I__11440 (
            .O(N__49147),
            .I(N__48825));
    ClkMux I__11439 (
            .O(N__49146),
            .I(N__48825));
    ClkMux I__11438 (
            .O(N__49145),
            .I(N__48825));
    ClkMux I__11437 (
            .O(N__49144),
            .I(N__48825));
    ClkMux I__11436 (
            .O(N__49143),
            .I(N__48825));
    ClkMux I__11435 (
            .O(N__49142),
            .I(N__48825));
    ClkMux I__11434 (
            .O(N__49141),
            .I(N__48825));
    ClkMux I__11433 (
            .O(N__49140),
            .I(N__48825));
    ClkMux I__11432 (
            .O(N__49139),
            .I(N__48825));
    ClkMux I__11431 (
            .O(N__49138),
            .I(N__48825));
    ClkMux I__11430 (
            .O(N__49137),
            .I(N__48825));
    ClkMux I__11429 (
            .O(N__49136),
            .I(N__48825));
    ClkMux I__11428 (
            .O(N__49135),
            .I(N__48825));
    ClkMux I__11427 (
            .O(N__49134),
            .I(N__48825));
    ClkMux I__11426 (
            .O(N__49133),
            .I(N__48825));
    ClkMux I__11425 (
            .O(N__49132),
            .I(N__48825));
    ClkMux I__11424 (
            .O(N__49131),
            .I(N__48825));
    ClkMux I__11423 (
            .O(N__49130),
            .I(N__48825));
    ClkMux I__11422 (
            .O(N__49129),
            .I(N__48825));
    ClkMux I__11421 (
            .O(N__49128),
            .I(N__48825));
    ClkMux I__11420 (
            .O(N__49127),
            .I(N__48825));
    ClkMux I__11419 (
            .O(N__49126),
            .I(N__48825));
    ClkMux I__11418 (
            .O(N__49125),
            .I(N__48825));
    ClkMux I__11417 (
            .O(N__49124),
            .I(N__48825));
    ClkMux I__11416 (
            .O(N__49123),
            .I(N__48825));
    ClkMux I__11415 (
            .O(N__49122),
            .I(N__48825));
    ClkMux I__11414 (
            .O(N__49121),
            .I(N__48825));
    ClkMux I__11413 (
            .O(N__49120),
            .I(N__48825));
    ClkMux I__11412 (
            .O(N__49119),
            .I(N__48825));
    ClkMux I__11411 (
            .O(N__49118),
            .I(N__48825));
    ClkMux I__11410 (
            .O(N__49117),
            .I(N__48825));
    ClkMux I__11409 (
            .O(N__49116),
            .I(N__48825));
    ClkMux I__11408 (
            .O(N__49115),
            .I(N__48825));
    ClkMux I__11407 (
            .O(N__49114),
            .I(N__48825));
    ClkMux I__11406 (
            .O(N__49113),
            .I(N__48825));
    ClkMux I__11405 (
            .O(N__49112),
            .I(N__48825));
    ClkMux I__11404 (
            .O(N__49111),
            .I(N__48825));
    ClkMux I__11403 (
            .O(N__49110),
            .I(N__48825));
    GlobalMux I__11402 (
            .O(N__48825),
            .I(clk_100mhz_0));
    CEMux I__11401 (
            .O(N__48822),
            .I(N__48816));
    CEMux I__11400 (
            .O(N__48821),
            .I(N__48808));
    CEMux I__11399 (
            .O(N__48820),
            .I(N__48798));
    CEMux I__11398 (
            .O(N__48819),
            .I(N__48795));
    LocalMux I__11397 (
            .O(N__48816),
            .I(N__48792));
    InMux I__11396 (
            .O(N__48815),
            .I(N__48783));
    InMux I__11395 (
            .O(N__48814),
            .I(N__48783));
    InMux I__11394 (
            .O(N__48813),
            .I(N__48783));
    InMux I__11393 (
            .O(N__48812),
            .I(N__48783));
    CEMux I__11392 (
            .O(N__48811),
            .I(N__48780));
    LocalMux I__11391 (
            .O(N__48808),
            .I(N__48777));
    InMux I__11390 (
            .O(N__48807),
            .I(N__48770));
    InMux I__11389 (
            .O(N__48806),
            .I(N__48770));
    InMux I__11388 (
            .O(N__48805),
            .I(N__48770));
    CEMux I__11387 (
            .O(N__48804),
            .I(N__48767));
    CEMux I__11386 (
            .O(N__48803),
            .I(N__48764));
    CEMux I__11385 (
            .O(N__48802),
            .I(N__48742));
    CEMux I__11384 (
            .O(N__48801),
            .I(N__48739));
    LocalMux I__11383 (
            .O(N__48798),
            .I(N__48736));
    LocalMux I__11382 (
            .O(N__48795),
            .I(N__48733));
    Span4Mux_h I__11381 (
            .O(N__48792),
            .I(N__48730));
    LocalMux I__11380 (
            .O(N__48783),
            .I(N__48727));
    LocalMux I__11379 (
            .O(N__48780),
            .I(N__48722));
    Span4Mux_v I__11378 (
            .O(N__48777),
            .I(N__48722));
    LocalMux I__11377 (
            .O(N__48770),
            .I(N__48717));
    LocalMux I__11376 (
            .O(N__48767),
            .I(N__48717));
    LocalMux I__11375 (
            .O(N__48764),
            .I(N__48714));
    InMux I__11374 (
            .O(N__48763),
            .I(N__48705));
    InMux I__11373 (
            .O(N__48762),
            .I(N__48705));
    InMux I__11372 (
            .O(N__48761),
            .I(N__48705));
    InMux I__11371 (
            .O(N__48760),
            .I(N__48705));
    InMux I__11370 (
            .O(N__48759),
            .I(N__48696));
    InMux I__11369 (
            .O(N__48758),
            .I(N__48696));
    InMux I__11368 (
            .O(N__48757),
            .I(N__48696));
    InMux I__11367 (
            .O(N__48756),
            .I(N__48696));
    InMux I__11366 (
            .O(N__48755),
            .I(N__48689));
    InMux I__11365 (
            .O(N__48754),
            .I(N__48689));
    InMux I__11364 (
            .O(N__48753),
            .I(N__48689));
    InMux I__11363 (
            .O(N__48752),
            .I(N__48680));
    InMux I__11362 (
            .O(N__48751),
            .I(N__48680));
    InMux I__11361 (
            .O(N__48750),
            .I(N__48680));
    InMux I__11360 (
            .O(N__48749),
            .I(N__48680));
    InMux I__11359 (
            .O(N__48748),
            .I(N__48671));
    InMux I__11358 (
            .O(N__48747),
            .I(N__48671));
    InMux I__11357 (
            .O(N__48746),
            .I(N__48671));
    InMux I__11356 (
            .O(N__48745),
            .I(N__48671));
    LocalMux I__11355 (
            .O(N__48742),
            .I(N__48663));
    LocalMux I__11354 (
            .O(N__48739),
            .I(N__48660));
    Span4Mux_v I__11353 (
            .O(N__48736),
            .I(N__48655));
    Span4Mux_v I__11352 (
            .O(N__48733),
            .I(N__48655));
    Span4Mux_v I__11351 (
            .O(N__48730),
            .I(N__48652));
    Span4Mux_v I__11350 (
            .O(N__48727),
            .I(N__48645));
    Span4Mux_v I__11349 (
            .O(N__48722),
            .I(N__48645));
    Span4Mux_v I__11348 (
            .O(N__48717),
            .I(N__48645));
    Span4Mux_v I__11347 (
            .O(N__48714),
            .I(N__48638));
    LocalMux I__11346 (
            .O(N__48705),
            .I(N__48638));
    LocalMux I__11345 (
            .O(N__48696),
            .I(N__48638));
    LocalMux I__11344 (
            .O(N__48689),
            .I(N__48631));
    LocalMux I__11343 (
            .O(N__48680),
            .I(N__48631));
    LocalMux I__11342 (
            .O(N__48671),
            .I(N__48631));
    InMux I__11341 (
            .O(N__48670),
            .I(N__48622));
    InMux I__11340 (
            .O(N__48669),
            .I(N__48622));
    InMux I__11339 (
            .O(N__48668),
            .I(N__48622));
    InMux I__11338 (
            .O(N__48667),
            .I(N__48622));
    InMux I__11337 (
            .O(N__48666),
            .I(N__48619));
    Sp12to4 I__11336 (
            .O(N__48663),
            .I(N__48616));
    Span4Mux_v I__11335 (
            .O(N__48660),
            .I(N__48611));
    Span4Mux_v I__11334 (
            .O(N__48655),
            .I(N__48611));
    Span4Mux_h I__11333 (
            .O(N__48652),
            .I(N__48602));
    Span4Mux_h I__11332 (
            .O(N__48645),
            .I(N__48602));
    Span4Mux_v I__11331 (
            .O(N__48638),
            .I(N__48602));
    Span4Mux_v I__11330 (
            .O(N__48631),
            .I(N__48602));
    LocalMux I__11329 (
            .O(N__48622),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    LocalMux I__11328 (
            .O(N__48619),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv12 I__11327 (
            .O(N__48616),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11326 (
            .O(N__48611),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11325 (
            .O(N__48602),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__11324 (
            .O(N__48591),
            .I(N__48580));
    InMux I__11323 (
            .O(N__48590),
            .I(N__48577));
    InMux I__11322 (
            .O(N__48589),
            .I(N__48574));
    InMux I__11321 (
            .O(N__48588),
            .I(N__48571));
    InMux I__11320 (
            .O(N__48587),
            .I(N__48568));
    InMux I__11319 (
            .O(N__48586),
            .I(N__48565));
    InMux I__11318 (
            .O(N__48585),
            .I(N__48562));
    InMux I__11317 (
            .O(N__48584),
            .I(N__48559));
    InMux I__11316 (
            .O(N__48583),
            .I(N__48556));
    LocalMux I__11315 (
            .O(N__48580),
            .I(N__48553));
    LocalMux I__11314 (
            .O(N__48577),
            .I(N__48550));
    LocalMux I__11313 (
            .O(N__48574),
            .I(N__48547));
    LocalMux I__11312 (
            .O(N__48571),
            .I(N__48501));
    LocalMux I__11311 (
            .O(N__48568),
            .I(N__48489));
    LocalMux I__11310 (
            .O(N__48565),
            .I(N__48450));
    LocalMux I__11309 (
            .O(N__48562),
            .I(N__48438));
    LocalMux I__11308 (
            .O(N__48559),
            .I(N__48423));
    LocalMux I__11307 (
            .O(N__48556),
            .I(N__48409));
    Glb2LocalMux I__11306 (
            .O(N__48553),
            .I(N__48096));
    Glb2LocalMux I__11305 (
            .O(N__48550),
            .I(N__48096));
    Glb2LocalMux I__11304 (
            .O(N__48547),
            .I(N__48096));
    SRMux I__11303 (
            .O(N__48546),
            .I(N__48096));
    SRMux I__11302 (
            .O(N__48545),
            .I(N__48096));
    SRMux I__11301 (
            .O(N__48544),
            .I(N__48096));
    SRMux I__11300 (
            .O(N__48543),
            .I(N__48096));
    SRMux I__11299 (
            .O(N__48542),
            .I(N__48096));
    SRMux I__11298 (
            .O(N__48541),
            .I(N__48096));
    SRMux I__11297 (
            .O(N__48540),
            .I(N__48096));
    SRMux I__11296 (
            .O(N__48539),
            .I(N__48096));
    SRMux I__11295 (
            .O(N__48538),
            .I(N__48096));
    SRMux I__11294 (
            .O(N__48537),
            .I(N__48096));
    SRMux I__11293 (
            .O(N__48536),
            .I(N__48096));
    SRMux I__11292 (
            .O(N__48535),
            .I(N__48096));
    SRMux I__11291 (
            .O(N__48534),
            .I(N__48096));
    SRMux I__11290 (
            .O(N__48533),
            .I(N__48096));
    SRMux I__11289 (
            .O(N__48532),
            .I(N__48096));
    SRMux I__11288 (
            .O(N__48531),
            .I(N__48096));
    SRMux I__11287 (
            .O(N__48530),
            .I(N__48096));
    SRMux I__11286 (
            .O(N__48529),
            .I(N__48096));
    SRMux I__11285 (
            .O(N__48528),
            .I(N__48096));
    SRMux I__11284 (
            .O(N__48527),
            .I(N__48096));
    SRMux I__11283 (
            .O(N__48526),
            .I(N__48096));
    SRMux I__11282 (
            .O(N__48525),
            .I(N__48096));
    SRMux I__11281 (
            .O(N__48524),
            .I(N__48096));
    SRMux I__11280 (
            .O(N__48523),
            .I(N__48096));
    SRMux I__11279 (
            .O(N__48522),
            .I(N__48096));
    SRMux I__11278 (
            .O(N__48521),
            .I(N__48096));
    SRMux I__11277 (
            .O(N__48520),
            .I(N__48096));
    SRMux I__11276 (
            .O(N__48519),
            .I(N__48096));
    SRMux I__11275 (
            .O(N__48518),
            .I(N__48096));
    SRMux I__11274 (
            .O(N__48517),
            .I(N__48096));
    SRMux I__11273 (
            .O(N__48516),
            .I(N__48096));
    SRMux I__11272 (
            .O(N__48515),
            .I(N__48096));
    SRMux I__11271 (
            .O(N__48514),
            .I(N__48096));
    SRMux I__11270 (
            .O(N__48513),
            .I(N__48096));
    SRMux I__11269 (
            .O(N__48512),
            .I(N__48096));
    SRMux I__11268 (
            .O(N__48511),
            .I(N__48096));
    SRMux I__11267 (
            .O(N__48510),
            .I(N__48096));
    SRMux I__11266 (
            .O(N__48509),
            .I(N__48096));
    SRMux I__11265 (
            .O(N__48508),
            .I(N__48096));
    SRMux I__11264 (
            .O(N__48507),
            .I(N__48096));
    SRMux I__11263 (
            .O(N__48506),
            .I(N__48096));
    SRMux I__11262 (
            .O(N__48505),
            .I(N__48096));
    SRMux I__11261 (
            .O(N__48504),
            .I(N__48096));
    Glb2LocalMux I__11260 (
            .O(N__48501),
            .I(N__48096));
    SRMux I__11259 (
            .O(N__48500),
            .I(N__48096));
    SRMux I__11258 (
            .O(N__48499),
            .I(N__48096));
    SRMux I__11257 (
            .O(N__48498),
            .I(N__48096));
    SRMux I__11256 (
            .O(N__48497),
            .I(N__48096));
    SRMux I__11255 (
            .O(N__48496),
            .I(N__48096));
    SRMux I__11254 (
            .O(N__48495),
            .I(N__48096));
    SRMux I__11253 (
            .O(N__48494),
            .I(N__48096));
    SRMux I__11252 (
            .O(N__48493),
            .I(N__48096));
    SRMux I__11251 (
            .O(N__48492),
            .I(N__48096));
    Glb2LocalMux I__11250 (
            .O(N__48489),
            .I(N__48096));
    SRMux I__11249 (
            .O(N__48488),
            .I(N__48096));
    SRMux I__11248 (
            .O(N__48487),
            .I(N__48096));
    SRMux I__11247 (
            .O(N__48486),
            .I(N__48096));
    SRMux I__11246 (
            .O(N__48485),
            .I(N__48096));
    SRMux I__11245 (
            .O(N__48484),
            .I(N__48096));
    SRMux I__11244 (
            .O(N__48483),
            .I(N__48096));
    SRMux I__11243 (
            .O(N__48482),
            .I(N__48096));
    SRMux I__11242 (
            .O(N__48481),
            .I(N__48096));
    SRMux I__11241 (
            .O(N__48480),
            .I(N__48096));
    SRMux I__11240 (
            .O(N__48479),
            .I(N__48096));
    SRMux I__11239 (
            .O(N__48478),
            .I(N__48096));
    SRMux I__11238 (
            .O(N__48477),
            .I(N__48096));
    SRMux I__11237 (
            .O(N__48476),
            .I(N__48096));
    SRMux I__11236 (
            .O(N__48475),
            .I(N__48096));
    SRMux I__11235 (
            .O(N__48474),
            .I(N__48096));
    SRMux I__11234 (
            .O(N__48473),
            .I(N__48096));
    SRMux I__11233 (
            .O(N__48472),
            .I(N__48096));
    SRMux I__11232 (
            .O(N__48471),
            .I(N__48096));
    SRMux I__11231 (
            .O(N__48470),
            .I(N__48096));
    SRMux I__11230 (
            .O(N__48469),
            .I(N__48096));
    SRMux I__11229 (
            .O(N__48468),
            .I(N__48096));
    SRMux I__11228 (
            .O(N__48467),
            .I(N__48096));
    SRMux I__11227 (
            .O(N__48466),
            .I(N__48096));
    SRMux I__11226 (
            .O(N__48465),
            .I(N__48096));
    SRMux I__11225 (
            .O(N__48464),
            .I(N__48096));
    SRMux I__11224 (
            .O(N__48463),
            .I(N__48096));
    SRMux I__11223 (
            .O(N__48462),
            .I(N__48096));
    SRMux I__11222 (
            .O(N__48461),
            .I(N__48096));
    SRMux I__11221 (
            .O(N__48460),
            .I(N__48096));
    SRMux I__11220 (
            .O(N__48459),
            .I(N__48096));
    SRMux I__11219 (
            .O(N__48458),
            .I(N__48096));
    SRMux I__11218 (
            .O(N__48457),
            .I(N__48096));
    SRMux I__11217 (
            .O(N__48456),
            .I(N__48096));
    SRMux I__11216 (
            .O(N__48455),
            .I(N__48096));
    SRMux I__11215 (
            .O(N__48454),
            .I(N__48096));
    SRMux I__11214 (
            .O(N__48453),
            .I(N__48096));
    Glb2LocalMux I__11213 (
            .O(N__48450),
            .I(N__48096));
    SRMux I__11212 (
            .O(N__48449),
            .I(N__48096));
    SRMux I__11211 (
            .O(N__48448),
            .I(N__48096));
    SRMux I__11210 (
            .O(N__48447),
            .I(N__48096));
    SRMux I__11209 (
            .O(N__48446),
            .I(N__48096));
    SRMux I__11208 (
            .O(N__48445),
            .I(N__48096));
    SRMux I__11207 (
            .O(N__48444),
            .I(N__48096));
    SRMux I__11206 (
            .O(N__48443),
            .I(N__48096));
    SRMux I__11205 (
            .O(N__48442),
            .I(N__48096));
    SRMux I__11204 (
            .O(N__48441),
            .I(N__48096));
    Glb2LocalMux I__11203 (
            .O(N__48438),
            .I(N__48096));
    SRMux I__11202 (
            .O(N__48437),
            .I(N__48096));
    SRMux I__11201 (
            .O(N__48436),
            .I(N__48096));
    SRMux I__11200 (
            .O(N__48435),
            .I(N__48096));
    SRMux I__11199 (
            .O(N__48434),
            .I(N__48096));
    SRMux I__11198 (
            .O(N__48433),
            .I(N__48096));
    SRMux I__11197 (
            .O(N__48432),
            .I(N__48096));
    SRMux I__11196 (
            .O(N__48431),
            .I(N__48096));
    SRMux I__11195 (
            .O(N__48430),
            .I(N__48096));
    SRMux I__11194 (
            .O(N__48429),
            .I(N__48096));
    SRMux I__11193 (
            .O(N__48428),
            .I(N__48096));
    SRMux I__11192 (
            .O(N__48427),
            .I(N__48096));
    SRMux I__11191 (
            .O(N__48426),
            .I(N__48096));
    Glb2LocalMux I__11190 (
            .O(N__48423),
            .I(N__48096));
    SRMux I__11189 (
            .O(N__48422),
            .I(N__48096));
    SRMux I__11188 (
            .O(N__48421),
            .I(N__48096));
    SRMux I__11187 (
            .O(N__48420),
            .I(N__48096));
    SRMux I__11186 (
            .O(N__48419),
            .I(N__48096));
    SRMux I__11185 (
            .O(N__48418),
            .I(N__48096));
    SRMux I__11184 (
            .O(N__48417),
            .I(N__48096));
    SRMux I__11183 (
            .O(N__48416),
            .I(N__48096));
    SRMux I__11182 (
            .O(N__48415),
            .I(N__48096));
    SRMux I__11181 (
            .O(N__48414),
            .I(N__48096));
    SRMux I__11180 (
            .O(N__48413),
            .I(N__48096));
    SRMux I__11179 (
            .O(N__48412),
            .I(N__48096));
    Glb2LocalMux I__11178 (
            .O(N__48409),
            .I(N__48096));
    SRMux I__11177 (
            .O(N__48408),
            .I(N__48096));
    SRMux I__11176 (
            .O(N__48407),
            .I(N__48096));
    SRMux I__11175 (
            .O(N__48406),
            .I(N__48096));
    SRMux I__11174 (
            .O(N__48405),
            .I(N__48096));
    SRMux I__11173 (
            .O(N__48404),
            .I(N__48096));
    SRMux I__11172 (
            .O(N__48403),
            .I(N__48096));
    SRMux I__11171 (
            .O(N__48402),
            .I(N__48096));
    SRMux I__11170 (
            .O(N__48401),
            .I(N__48096));
    SRMux I__11169 (
            .O(N__48400),
            .I(N__48096));
    SRMux I__11168 (
            .O(N__48399),
            .I(N__48096));
    SRMux I__11167 (
            .O(N__48398),
            .I(N__48096));
    SRMux I__11166 (
            .O(N__48397),
            .I(N__48096));
    SRMux I__11165 (
            .O(N__48396),
            .I(N__48096));
    SRMux I__11164 (
            .O(N__48395),
            .I(N__48096));
    SRMux I__11163 (
            .O(N__48394),
            .I(N__48096));
    SRMux I__11162 (
            .O(N__48393),
            .I(N__48096));
    SRMux I__11161 (
            .O(N__48392),
            .I(N__48096));
    SRMux I__11160 (
            .O(N__48391),
            .I(N__48096));
    GlobalMux I__11159 (
            .O(N__48096),
            .I(N__48093));
    gio2CtrlBuf I__11158 (
            .O(N__48093),
            .I(red_c_g));
    InMux I__11157 (
            .O(N__48090),
            .I(N__48052));
    InMux I__11156 (
            .O(N__48089),
            .I(N__48052));
    InMux I__11155 (
            .O(N__48088),
            .I(N__48052));
    InMux I__11154 (
            .O(N__48087),
            .I(N__48052));
    InMux I__11153 (
            .O(N__48086),
            .I(N__48043));
    InMux I__11152 (
            .O(N__48085),
            .I(N__48043));
    InMux I__11151 (
            .O(N__48084),
            .I(N__48043));
    InMux I__11150 (
            .O(N__48083),
            .I(N__48043));
    InMux I__11149 (
            .O(N__48082),
            .I(N__48038));
    InMux I__11148 (
            .O(N__48081),
            .I(N__48038));
    InMux I__11147 (
            .O(N__48080),
            .I(N__48029));
    InMux I__11146 (
            .O(N__48079),
            .I(N__48029));
    InMux I__11145 (
            .O(N__48078),
            .I(N__48029));
    InMux I__11144 (
            .O(N__48077),
            .I(N__48029));
    InMux I__11143 (
            .O(N__48076),
            .I(N__48020));
    InMux I__11142 (
            .O(N__48075),
            .I(N__48020));
    InMux I__11141 (
            .O(N__48074),
            .I(N__48020));
    InMux I__11140 (
            .O(N__48073),
            .I(N__48020));
    InMux I__11139 (
            .O(N__48072),
            .I(N__48011));
    InMux I__11138 (
            .O(N__48071),
            .I(N__48011));
    InMux I__11137 (
            .O(N__48070),
            .I(N__48011));
    InMux I__11136 (
            .O(N__48069),
            .I(N__48011));
    InMux I__11135 (
            .O(N__48068),
            .I(N__48002));
    InMux I__11134 (
            .O(N__48067),
            .I(N__48002));
    InMux I__11133 (
            .O(N__48066),
            .I(N__48002));
    InMux I__11132 (
            .O(N__48065),
            .I(N__48002));
    InMux I__11131 (
            .O(N__48064),
            .I(N__47993));
    InMux I__11130 (
            .O(N__48063),
            .I(N__47993));
    InMux I__11129 (
            .O(N__48062),
            .I(N__47993));
    InMux I__11128 (
            .O(N__48061),
            .I(N__47993));
    LocalMux I__11127 (
            .O(N__48052),
            .I(N__47990));
    LocalMux I__11126 (
            .O(N__48043),
            .I(N__47987));
    LocalMux I__11125 (
            .O(N__48038),
            .I(N__47974));
    LocalMux I__11124 (
            .O(N__48029),
            .I(N__47974));
    LocalMux I__11123 (
            .O(N__48020),
            .I(N__47974));
    LocalMux I__11122 (
            .O(N__48011),
            .I(N__47974));
    LocalMux I__11121 (
            .O(N__48002),
            .I(N__47974));
    LocalMux I__11120 (
            .O(N__47993),
            .I(N__47974));
    Span4Mux_h I__11119 (
            .O(N__47990),
            .I(N__47971));
    Span4Mux_v I__11118 (
            .O(N__47987),
            .I(N__47966));
    Span4Mux_v I__11117 (
            .O(N__47974),
            .I(N__47966));
    Odrv4 I__11116 (
            .O(N__47971),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__11115 (
            .O(N__47966),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__11114 (
            .O(N__47961),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__11113 (
            .O(N__47958),
            .I(N__47954));
    InMux I__11112 (
            .O(N__47957),
            .I(N__47951));
    LocalMux I__11111 (
            .O(N__47954),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__11110 (
            .O(N__47951),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__11109 (
            .O(N__47946),
            .I(N__47941));
    CEMux I__11108 (
            .O(N__47945),
            .I(N__47938));
    CEMux I__11107 (
            .O(N__47944),
            .I(N__47935));
    LocalMux I__11106 (
            .O(N__47941),
            .I(N__47929));
    LocalMux I__11105 (
            .O(N__47938),
            .I(N__47929));
    LocalMux I__11104 (
            .O(N__47935),
            .I(N__47926));
    CEMux I__11103 (
            .O(N__47934),
            .I(N__47923));
    Span4Mux_v I__11102 (
            .O(N__47929),
            .I(N__47920));
    Span4Mux_v I__11101 (
            .O(N__47926),
            .I(N__47915));
    LocalMux I__11100 (
            .O(N__47923),
            .I(N__47915));
    Span4Mux_h I__11099 (
            .O(N__47920),
            .I(N__47910));
    Span4Mux_h I__11098 (
            .O(N__47915),
            .I(N__47910));
    Odrv4 I__11097 (
            .O(N__47910),
            .I(\delay_measurement_inst.delay_tr_timer.N_396_i ));
    CascadeMux I__11096 (
            .O(N__47907),
            .I(N__47904));
    InMux I__11095 (
            .O(N__47904),
            .I(N__47901));
    LocalMux I__11094 (
            .O(N__47901),
            .I(N__47898));
    Span12Mux_v I__11093 (
            .O(N__47898),
            .I(N__47894));
    InMux I__11092 (
            .O(N__47897),
            .I(N__47891));
    Odrv12 I__11091 (
            .O(N__47894),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__11090 (
            .O(N__47891),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__11089 (
            .O(N__47886),
            .I(N__47882));
    InMux I__11088 (
            .O(N__47885),
            .I(N__47878));
    LocalMux I__11087 (
            .O(N__47882),
            .I(N__47875));
    InMux I__11086 (
            .O(N__47881),
            .I(N__47872));
    LocalMux I__11085 (
            .O(N__47878),
            .I(N__47868));
    Span4Mux_v I__11084 (
            .O(N__47875),
            .I(N__47863));
    LocalMux I__11083 (
            .O(N__47872),
            .I(N__47863));
    InMux I__11082 (
            .O(N__47871),
            .I(N__47860));
    Span4Mux_h I__11081 (
            .O(N__47868),
            .I(N__47857));
    Span4Mux_h I__11080 (
            .O(N__47863),
            .I(N__47854));
    LocalMux I__11079 (
            .O(N__47860),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    Odrv4 I__11078 (
            .O(N__47857),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    Odrv4 I__11077 (
            .O(N__47854),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    InMux I__11076 (
            .O(N__47847),
            .I(N__47843));
    InMux I__11075 (
            .O(N__47846),
            .I(N__47838));
    LocalMux I__11074 (
            .O(N__47843),
            .I(N__47835));
    InMux I__11073 (
            .O(N__47842),
            .I(N__47832));
    InMux I__11072 (
            .O(N__47841),
            .I(N__47829));
    LocalMux I__11071 (
            .O(N__47838),
            .I(N__47823));
    Span4Mux_v I__11070 (
            .O(N__47835),
            .I(N__47819));
    LocalMux I__11069 (
            .O(N__47832),
            .I(N__47814));
    LocalMux I__11068 (
            .O(N__47829),
            .I(N__47814));
    InMux I__11067 (
            .O(N__47828),
            .I(N__47807));
    InMux I__11066 (
            .O(N__47827),
            .I(N__47807));
    InMux I__11065 (
            .O(N__47826),
            .I(N__47807));
    Span4Mux_v I__11064 (
            .O(N__47823),
            .I(N__47804));
    InMux I__11063 (
            .O(N__47822),
            .I(N__47801));
    Span4Mux_h I__11062 (
            .O(N__47819),
            .I(N__47796));
    Span4Mux_v I__11061 (
            .O(N__47814),
            .I(N__47796));
    LocalMux I__11060 (
            .O(N__47807),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    Odrv4 I__11059 (
            .O(N__47804),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    LocalMux I__11058 (
            .O(N__47801),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    Odrv4 I__11057 (
            .O(N__47796),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    CascadeMux I__11056 (
            .O(N__47787),
            .I(elapsed_time_ns_1_RNII6NQL1_0_1_cascade_));
    InMux I__11055 (
            .O(N__47784),
            .I(N__47779));
    InMux I__11054 (
            .O(N__47783),
            .I(N__47776));
    InMux I__11053 (
            .O(N__47782),
            .I(N__47773));
    LocalMux I__11052 (
            .O(N__47779),
            .I(N__47770));
    LocalMux I__11051 (
            .O(N__47776),
            .I(N__47767));
    LocalMux I__11050 (
            .O(N__47773),
            .I(N__47763));
    Span4Mux_h I__11049 (
            .O(N__47770),
            .I(N__47760));
    Sp12to4 I__11048 (
            .O(N__47767),
            .I(N__47757));
    InMux I__11047 (
            .O(N__47766),
            .I(N__47754));
    Span4Mux_h I__11046 (
            .O(N__47763),
            .I(N__47751));
    Odrv4 I__11045 (
            .O(N__47760),
            .I(elapsed_time_ns_1_RNIBA65M1_0_19));
    Odrv12 I__11044 (
            .O(N__47757),
            .I(elapsed_time_ns_1_RNIBA65M1_0_19));
    LocalMux I__11043 (
            .O(N__47754),
            .I(elapsed_time_ns_1_RNIBA65M1_0_19));
    Odrv4 I__11042 (
            .O(N__47751),
            .I(elapsed_time_ns_1_RNIBA65M1_0_19));
    InMux I__11041 (
            .O(N__47742),
            .I(N__47739));
    LocalMux I__11040 (
            .O(N__47739),
            .I(N__47736));
    Span4Mux_v I__11039 (
            .O(N__47736),
            .I(N__47732));
    InMux I__11038 (
            .O(N__47735),
            .I(N__47729));
    Span4Mux_h I__11037 (
            .O(N__47732),
            .I(N__47723));
    LocalMux I__11036 (
            .O(N__47729),
            .I(N__47723));
    InMux I__11035 (
            .O(N__47728),
            .I(N__47720));
    Odrv4 I__11034 (
            .O(N__47723),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    LocalMux I__11033 (
            .O(N__47720),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__11032 (
            .O(N__47715),
            .I(N__47712));
    LocalMux I__11031 (
            .O(N__47712),
            .I(N__47709));
    Span4Mux_h I__11030 (
            .O(N__47709),
            .I(N__47706));
    Odrv4 I__11029 (
            .O(N__47706),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ));
    InMux I__11028 (
            .O(N__47703),
            .I(N__47695));
    InMux I__11027 (
            .O(N__47702),
            .I(N__47692));
    CascadeMux I__11026 (
            .O(N__47701),
            .I(N__47687));
    InMux I__11025 (
            .O(N__47700),
            .I(N__47684));
    InMux I__11024 (
            .O(N__47699),
            .I(N__47681));
    InMux I__11023 (
            .O(N__47698),
            .I(N__47678));
    LocalMux I__11022 (
            .O(N__47695),
            .I(N__47672));
    LocalMux I__11021 (
            .O(N__47692),
            .I(N__47672));
    InMux I__11020 (
            .O(N__47691),
            .I(N__47669));
    InMux I__11019 (
            .O(N__47690),
            .I(N__47663));
    InMux I__11018 (
            .O(N__47687),
            .I(N__47663));
    LocalMux I__11017 (
            .O(N__47684),
            .I(N__47659));
    LocalMux I__11016 (
            .O(N__47681),
            .I(N__47656));
    LocalMux I__11015 (
            .O(N__47678),
            .I(N__47653));
    InMux I__11014 (
            .O(N__47677),
            .I(N__47650));
    Span4Mux_v I__11013 (
            .O(N__47672),
            .I(N__47645));
    LocalMux I__11012 (
            .O(N__47669),
            .I(N__47645));
    InMux I__11011 (
            .O(N__47668),
            .I(N__47641));
    LocalMux I__11010 (
            .O(N__47663),
            .I(N__47638));
    InMux I__11009 (
            .O(N__47662),
            .I(N__47635));
    Span4Mux_v I__11008 (
            .O(N__47659),
            .I(N__47627));
    Span4Mux_v I__11007 (
            .O(N__47656),
            .I(N__47619));
    Span4Mux_v I__11006 (
            .O(N__47653),
            .I(N__47619));
    LocalMux I__11005 (
            .O(N__47650),
            .I(N__47619));
    Span4Mux_h I__11004 (
            .O(N__47645),
            .I(N__47616));
    CascadeMux I__11003 (
            .O(N__47644),
            .I(N__47612));
    LocalMux I__11002 (
            .O(N__47641),
            .I(N__47605));
    Span4Mux_h I__11001 (
            .O(N__47638),
            .I(N__47605));
    LocalMux I__11000 (
            .O(N__47635),
            .I(N__47602));
    InMux I__10999 (
            .O(N__47634),
            .I(N__47597));
    InMux I__10998 (
            .O(N__47633),
            .I(N__47597));
    InMux I__10997 (
            .O(N__47632),
            .I(N__47590));
    InMux I__10996 (
            .O(N__47631),
            .I(N__47590));
    InMux I__10995 (
            .O(N__47630),
            .I(N__47590));
    Span4Mux_h I__10994 (
            .O(N__47627),
            .I(N__47587));
    InMux I__10993 (
            .O(N__47626),
            .I(N__47584));
    Span4Mux_h I__10992 (
            .O(N__47619),
            .I(N__47579));
    Span4Mux_v I__10991 (
            .O(N__47616),
            .I(N__47579));
    InMux I__10990 (
            .O(N__47615),
            .I(N__47576));
    InMux I__10989 (
            .O(N__47612),
            .I(N__47569));
    InMux I__10988 (
            .O(N__47611),
            .I(N__47569));
    InMux I__10987 (
            .O(N__47610),
            .I(N__47569));
    Span4Mux_h I__10986 (
            .O(N__47605),
            .I(N__47566));
    Span12Mux_v I__10985 (
            .O(N__47602),
            .I(N__47559));
    LocalMux I__10984 (
            .O(N__47597),
            .I(N__47559));
    LocalMux I__10983 (
            .O(N__47590),
            .I(N__47559));
    Odrv4 I__10982 (
            .O(N__47587),
            .I(\delay_measurement_inst.delay_tr9 ));
    LocalMux I__10981 (
            .O(N__47584),
            .I(\delay_measurement_inst.delay_tr9 ));
    Odrv4 I__10980 (
            .O(N__47579),
            .I(\delay_measurement_inst.delay_tr9 ));
    LocalMux I__10979 (
            .O(N__47576),
            .I(\delay_measurement_inst.delay_tr9 ));
    LocalMux I__10978 (
            .O(N__47569),
            .I(\delay_measurement_inst.delay_tr9 ));
    Odrv4 I__10977 (
            .O(N__47566),
            .I(\delay_measurement_inst.delay_tr9 ));
    Odrv12 I__10976 (
            .O(N__47559),
            .I(\delay_measurement_inst.delay_tr9 ));
    InMux I__10975 (
            .O(N__47544),
            .I(N__47541));
    LocalMux I__10974 (
            .O(N__47541),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1 ));
    CascadeMux I__10973 (
            .O(N__47538),
            .I(N__47534));
    InMux I__10972 (
            .O(N__47537),
            .I(N__47531));
    InMux I__10971 (
            .O(N__47534),
            .I(N__47528));
    LocalMux I__10970 (
            .O(N__47531),
            .I(N__47524));
    LocalMux I__10969 (
            .O(N__47528),
            .I(N__47521));
    InMux I__10968 (
            .O(N__47527),
            .I(N__47517));
    Span4Mux_v I__10967 (
            .O(N__47524),
            .I(N__47512));
    Span4Mux_v I__10966 (
            .O(N__47521),
            .I(N__47512));
    InMux I__10965 (
            .O(N__47520),
            .I(N__47509));
    LocalMux I__10964 (
            .O(N__47517),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    Odrv4 I__10963 (
            .O(N__47512),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    LocalMux I__10962 (
            .O(N__47509),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    InMux I__10961 (
            .O(N__47502),
            .I(N__47499));
    LocalMux I__10960 (
            .O(N__47499),
            .I(N__47496));
    Span12Mux_h I__10959 (
            .O(N__47496),
            .I(N__47493));
    Odrv12 I__10958 (
            .O(N__47493),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    InMux I__10957 (
            .O(N__47490),
            .I(N__47487));
    LocalMux I__10956 (
            .O(N__47487),
            .I(N__47484));
    Odrv12 I__10955 (
            .O(N__47484),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__10954 (
            .O(N__47481),
            .I(N__47478));
    InMux I__10953 (
            .O(N__47478),
            .I(N__47473));
    InMux I__10952 (
            .O(N__47477),
            .I(N__47470));
    InMux I__10951 (
            .O(N__47476),
            .I(N__47467));
    LocalMux I__10950 (
            .O(N__47473),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__10949 (
            .O(N__47470),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__10948 (
            .O(N__47467),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__10947 (
            .O(N__47460),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    CascadeMux I__10946 (
            .O(N__47457),
            .I(N__47454));
    InMux I__10945 (
            .O(N__47454),
            .I(N__47449));
    InMux I__10944 (
            .O(N__47453),
            .I(N__47446));
    InMux I__10943 (
            .O(N__47452),
            .I(N__47443));
    LocalMux I__10942 (
            .O(N__47449),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__10941 (
            .O(N__47446),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__10940 (
            .O(N__47443),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__10939 (
            .O(N__47436),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    CascadeMux I__10938 (
            .O(N__47433),
            .I(N__47430));
    InMux I__10937 (
            .O(N__47430),
            .I(N__47425));
    InMux I__10936 (
            .O(N__47429),
            .I(N__47422));
    InMux I__10935 (
            .O(N__47428),
            .I(N__47419));
    LocalMux I__10934 (
            .O(N__47425),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__10933 (
            .O(N__47422),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__10932 (
            .O(N__47419),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__10931 (
            .O(N__47412),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    CascadeMux I__10930 (
            .O(N__47409),
            .I(N__47406));
    InMux I__10929 (
            .O(N__47406),
            .I(N__47401));
    InMux I__10928 (
            .O(N__47405),
            .I(N__47398));
    InMux I__10927 (
            .O(N__47404),
            .I(N__47395));
    LocalMux I__10926 (
            .O(N__47401),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__10925 (
            .O(N__47398),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__10924 (
            .O(N__47395),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__10923 (
            .O(N__47388),
            .I(bfn_18_21_0_));
    CascadeMux I__10922 (
            .O(N__47385),
            .I(N__47382));
    InMux I__10921 (
            .O(N__47382),
            .I(N__47377));
    InMux I__10920 (
            .O(N__47381),
            .I(N__47374));
    InMux I__10919 (
            .O(N__47380),
            .I(N__47371));
    LocalMux I__10918 (
            .O(N__47377),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__10917 (
            .O(N__47374),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__10916 (
            .O(N__47371),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__10915 (
            .O(N__47364),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    CascadeMux I__10914 (
            .O(N__47361),
            .I(N__47358));
    InMux I__10913 (
            .O(N__47358),
            .I(N__47353));
    InMux I__10912 (
            .O(N__47357),
            .I(N__47350));
    InMux I__10911 (
            .O(N__47356),
            .I(N__47347));
    LocalMux I__10910 (
            .O(N__47353),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__10909 (
            .O(N__47350),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__10908 (
            .O(N__47347),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__10907 (
            .O(N__47340),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    CascadeMux I__10906 (
            .O(N__47337),
            .I(N__47334));
    InMux I__10905 (
            .O(N__47334),
            .I(N__47329));
    InMux I__10904 (
            .O(N__47333),
            .I(N__47326));
    InMux I__10903 (
            .O(N__47332),
            .I(N__47323));
    LocalMux I__10902 (
            .O(N__47329),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__10901 (
            .O(N__47326),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__10900 (
            .O(N__47323),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__10899 (
            .O(N__47316),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__10898 (
            .O(N__47313),
            .I(N__47309));
    InMux I__10897 (
            .O(N__47312),
            .I(N__47306));
    LocalMux I__10896 (
            .O(N__47309),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__10895 (
            .O(N__47306),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__10894 (
            .O(N__47301),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    CascadeMux I__10893 (
            .O(N__47298),
            .I(N__47295));
    InMux I__10892 (
            .O(N__47295),
            .I(N__47290));
    InMux I__10891 (
            .O(N__47294),
            .I(N__47287));
    InMux I__10890 (
            .O(N__47293),
            .I(N__47284));
    LocalMux I__10889 (
            .O(N__47290),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__10888 (
            .O(N__47287),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__10887 (
            .O(N__47284),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__10886 (
            .O(N__47277),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    CascadeMux I__10885 (
            .O(N__47274),
            .I(N__47271));
    InMux I__10884 (
            .O(N__47271),
            .I(N__47266));
    InMux I__10883 (
            .O(N__47270),
            .I(N__47263));
    InMux I__10882 (
            .O(N__47269),
            .I(N__47260));
    LocalMux I__10881 (
            .O(N__47266),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__10880 (
            .O(N__47263),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__10879 (
            .O(N__47260),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__10878 (
            .O(N__47253),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    CascadeMux I__10877 (
            .O(N__47250),
            .I(N__47247));
    InMux I__10876 (
            .O(N__47247),
            .I(N__47242));
    InMux I__10875 (
            .O(N__47246),
            .I(N__47239));
    InMux I__10874 (
            .O(N__47245),
            .I(N__47236));
    LocalMux I__10873 (
            .O(N__47242),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__10872 (
            .O(N__47239),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__10871 (
            .O(N__47236),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__10870 (
            .O(N__47229),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__10869 (
            .O(N__47226),
            .I(N__47223));
    InMux I__10868 (
            .O(N__47223),
            .I(N__47218));
    InMux I__10867 (
            .O(N__47222),
            .I(N__47215));
    InMux I__10866 (
            .O(N__47221),
            .I(N__47212));
    LocalMux I__10865 (
            .O(N__47218),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__10864 (
            .O(N__47215),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__10863 (
            .O(N__47212),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__10862 (
            .O(N__47205),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    CascadeMux I__10861 (
            .O(N__47202),
            .I(N__47199));
    InMux I__10860 (
            .O(N__47199),
            .I(N__47194));
    InMux I__10859 (
            .O(N__47198),
            .I(N__47191));
    InMux I__10858 (
            .O(N__47197),
            .I(N__47188));
    LocalMux I__10857 (
            .O(N__47194),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__10856 (
            .O(N__47191),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__10855 (
            .O(N__47188),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__10854 (
            .O(N__47181),
            .I(bfn_18_20_0_));
    CascadeMux I__10853 (
            .O(N__47178),
            .I(N__47175));
    InMux I__10852 (
            .O(N__47175),
            .I(N__47170));
    InMux I__10851 (
            .O(N__47174),
            .I(N__47167));
    InMux I__10850 (
            .O(N__47173),
            .I(N__47164));
    LocalMux I__10849 (
            .O(N__47170),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__10848 (
            .O(N__47167),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__10847 (
            .O(N__47164),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__10846 (
            .O(N__47157),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    CascadeMux I__10845 (
            .O(N__47154),
            .I(N__47151));
    InMux I__10844 (
            .O(N__47151),
            .I(N__47146));
    InMux I__10843 (
            .O(N__47150),
            .I(N__47143));
    InMux I__10842 (
            .O(N__47149),
            .I(N__47140));
    LocalMux I__10841 (
            .O(N__47146),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__10840 (
            .O(N__47143),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__10839 (
            .O(N__47140),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__10838 (
            .O(N__47133),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    CascadeMux I__10837 (
            .O(N__47130),
            .I(N__47127));
    InMux I__10836 (
            .O(N__47127),
            .I(N__47122));
    InMux I__10835 (
            .O(N__47126),
            .I(N__47119));
    InMux I__10834 (
            .O(N__47125),
            .I(N__47116));
    LocalMux I__10833 (
            .O(N__47122),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__10832 (
            .O(N__47119),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__10831 (
            .O(N__47116),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__10830 (
            .O(N__47109),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    CascadeMux I__10829 (
            .O(N__47106),
            .I(N__47103));
    InMux I__10828 (
            .O(N__47103),
            .I(N__47098));
    InMux I__10827 (
            .O(N__47102),
            .I(N__47095));
    InMux I__10826 (
            .O(N__47101),
            .I(N__47092));
    LocalMux I__10825 (
            .O(N__47098),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__10824 (
            .O(N__47095),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__10823 (
            .O(N__47092),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__10822 (
            .O(N__47085),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    CascadeMux I__10821 (
            .O(N__47082),
            .I(N__47079));
    InMux I__10820 (
            .O(N__47079),
            .I(N__47074));
    InMux I__10819 (
            .O(N__47078),
            .I(N__47071));
    InMux I__10818 (
            .O(N__47077),
            .I(N__47068));
    LocalMux I__10817 (
            .O(N__47074),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__10816 (
            .O(N__47071),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__10815 (
            .O(N__47068),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__10814 (
            .O(N__47061),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__10813 (
            .O(N__47058),
            .I(N__47055));
    InMux I__10812 (
            .O(N__47055),
            .I(N__47050));
    InMux I__10811 (
            .O(N__47054),
            .I(N__47047));
    InMux I__10810 (
            .O(N__47053),
            .I(N__47044));
    LocalMux I__10809 (
            .O(N__47050),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__10808 (
            .O(N__47047),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__10807 (
            .O(N__47044),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__10806 (
            .O(N__47037),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    CascadeMux I__10805 (
            .O(N__47034),
            .I(N__47031));
    InMux I__10804 (
            .O(N__47031),
            .I(N__47026));
    InMux I__10803 (
            .O(N__47030),
            .I(N__47023));
    InMux I__10802 (
            .O(N__47029),
            .I(N__47020));
    LocalMux I__10801 (
            .O(N__47026),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__10800 (
            .O(N__47023),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__10799 (
            .O(N__47020),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__10798 (
            .O(N__47013),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__10797 (
            .O(N__47010),
            .I(N__47007));
    InMux I__10796 (
            .O(N__47007),
            .I(N__47002));
    InMux I__10795 (
            .O(N__47006),
            .I(N__46999));
    InMux I__10794 (
            .O(N__47005),
            .I(N__46996));
    LocalMux I__10793 (
            .O(N__47002),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__10792 (
            .O(N__46999),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__10791 (
            .O(N__46996),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__10790 (
            .O(N__46989),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    CascadeMux I__10789 (
            .O(N__46986),
            .I(N__46983));
    InMux I__10788 (
            .O(N__46983),
            .I(N__46978));
    InMux I__10787 (
            .O(N__46982),
            .I(N__46975));
    InMux I__10786 (
            .O(N__46981),
            .I(N__46972));
    LocalMux I__10785 (
            .O(N__46978),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__10784 (
            .O(N__46975),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__10783 (
            .O(N__46972),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__10782 (
            .O(N__46965),
            .I(bfn_18_19_0_));
    CascadeMux I__10781 (
            .O(N__46962),
            .I(N__46959));
    InMux I__10780 (
            .O(N__46959),
            .I(N__46954));
    InMux I__10779 (
            .O(N__46958),
            .I(N__46951));
    InMux I__10778 (
            .O(N__46957),
            .I(N__46948));
    LocalMux I__10777 (
            .O(N__46954),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__10776 (
            .O(N__46951),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__10775 (
            .O(N__46948),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__10774 (
            .O(N__46941),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__10773 (
            .O(N__46938),
            .I(N__46935));
    InMux I__10772 (
            .O(N__46935),
            .I(N__46930));
    InMux I__10771 (
            .O(N__46934),
            .I(N__46927));
    InMux I__10770 (
            .O(N__46933),
            .I(N__46924));
    LocalMux I__10769 (
            .O(N__46930),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__10768 (
            .O(N__46927),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__10767 (
            .O(N__46924),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__10766 (
            .O(N__46917),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    CascadeMux I__10765 (
            .O(N__46914),
            .I(N__46911));
    InMux I__10764 (
            .O(N__46911),
            .I(N__46906));
    InMux I__10763 (
            .O(N__46910),
            .I(N__46903));
    InMux I__10762 (
            .O(N__46909),
            .I(N__46900));
    LocalMux I__10761 (
            .O(N__46906),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__10760 (
            .O(N__46903),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__10759 (
            .O(N__46900),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__10758 (
            .O(N__46893),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    CascadeMux I__10757 (
            .O(N__46890),
            .I(N__46887));
    InMux I__10756 (
            .O(N__46887),
            .I(N__46882));
    InMux I__10755 (
            .O(N__46886),
            .I(N__46879));
    InMux I__10754 (
            .O(N__46885),
            .I(N__46875));
    LocalMux I__10753 (
            .O(N__46882),
            .I(N__46869));
    LocalMux I__10752 (
            .O(N__46879),
            .I(N__46869));
    InMux I__10751 (
            .O(N__46878),
            .I(N__46864));
    LocalMux I__10750 (
            .O(N__46875),
            .I(N__46861));
    InMux I__10749 (
            .O(N__46874),
            .I(N__46857));
    Span4Mux_h I__10748 (
            .O(N__46869),
            .I(N__46854));
    InMux I__10747 (
            .O(N__46868),
            .I(N__46851));
    InMux I__10746 (
            .O(N__46867),
            .I(N__46848));
    LocalMux I__10745 (
            .O(N__46864),
            .I(N__46843));
    Span12Mux_v I__10744 (
            .O(N__46861),
            .I(N__46843));
    InMux I__10743 (
            .O(N__46860),
            .I(N__46840));
    LocalMux I__10742 (
            .O(N__46857),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    Odrv4 I__10741 (
            .O(N__46854),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__10740 (
            .O(N__46851),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__10739 (
            .O(N__46848),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    Odrv12 I__10738 (
            .O(N__46843),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__10737 (
            .O(N__46840),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    CascadeMux I__10736 (
            .O(N__46827),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_ ));
    InMux I__10735 (
            .O(N__46824),
            .I(N__46809));
    InMux I__10734 (
            .O(N__46823),
            .I(N__46804));
    InMux I__10733 (
            .O(N__46822),
            .I(N__46797));
    InMux I__10732 (
            .O(N__46821),
            .I(N__46797));
    InMux I__10731 (
            .O(N__46820),
            .I(N__46797));
    InMux I__10730 (
            .O(N__46819),
            .I(N__46794));
    InMux I__10729 (
            .O(N__46818),
            .I(N__46791));
    InMux I__10728 (
            .O(N__46817),
            .I(N__46784));
    InMux I__10727 (
            .O(N__46816),
            .I(N__46784));
    InMux I__10726 (
            .O(N__46815),
            .I(N__46784));
    InMux I__10725 (
            .O(N__46814),
            .I(N__46779));
    InMux I__10724 (
            .O(N__46813),
            .I(N__46779));
    InMux I__10723 (
            .O(N__46812),
            .I(N__46776));
    LocalMux I__10722 (
            .O(N__46809),
            .I(N__46773));
    CascadeMux I__10721 (
            .O(N__46808),
            .I(N__46769));
    CascadeMux I__10720 (
            .O(N__46807),
            .I(N__46761));
    LocalMux I__10719 (
            .O(N__46804),
            .I(N__46758));
    LocalMux I__10718 (
            .O(N__46797),
            .I(N__46753));
    LocalMux I__10717 (
            .O(N__46794),
            .I(N__46753));
    LocalMux I__10716 (
            .O(N__46791),
            .I(N__46745));
    LocalMux I__10715 (
            .O(N__46784),
            .I(N__46738));
    LocalMux I__10714 (
            .O(N__46779),
            .I(N__46738));
    LocalMux I__10713 (
            .O(N__46776),
            .I(N__46738));
    Span4Mux_v I__10712 (
            .O(N__46773),
            .I(N__46735));
    InMux I__10711 (
            .O(N__46772),
            .I(N__46728));
    InMux I__10710 (
            .O(N__46769),
            .I(N__46728));
    InMux I__10709 (
            .O(N__46768),
            .I(N__46728));
    InMux I__10708 (
            .O(N__46767),
            .I(N__46722));
    InMux I__10707 (
            .O(N__46766),
            .I(N__46722));
    InMux I__10706 (
            .O(N__46765),
            .I(N__46715));
    InMux I__10705 (
            .O(N__46764),
            .I(N__46715));
    InMux I__10704 (
            .O(N__46761),
            .I(N__46715));
    Span4Mux_h I__10703 (
            .O(N__46758),
            .I(N__46712));
    Span4Mux_v I__10702 (
            .O(N__46753),
            .I(N__46709));
    InMux I__10701 (
            .O(N__46752),
            .I(N__46698));
    InMux I__10700 (
            .O(N__46751),
            .I(N__46698));
    InMux I__10699 (
            .O(N__46750),
            .I(N__46698));
    InMux I__10698 (
            .O(N__46749),
            .I(N__46698));
    InMux I__10697 (
            .O(N__46748),
            .I(N__46698));
    Span4Mux_v I__10696 (
            .O(N__46745),
            .I(N__46689));
    Span4Mux_v I__10695 (
            .O(N__46738),
            .I(N__46689));
    Span4Mux_v I__10694 (
            .O(N__46735),
            .I(N__46689));
    LocalMux I__10693 (
            .O(N__46728),
            .I(N__46689));
    InMux I__10692 (
            .O(N__46727),
            .I(N__46686));
    LocalMux I__10691 (
            .O(N__46722),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__10690 (
            .O(N__46715),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv4 I__10689 (
            .O(N__46712),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv4 I__10688 (
            .O(N__46709),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__10687 (
            .O(N__46698),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv4 I__10686 (
            .O(N__46689),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    LocalMux I__10685 (
            .O(N__46686),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    CascadeMux I__10684 (
            .O(N__46671),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_ ));
    CascadeMux I__10683 (
            .O(N__46668),
            .I(N__46665));
    InMux I__10682 (
            .O(N__46665),
            .I(N__46662));
    LocalMux I__10681 (
            .O(N__46662),
            .I(N__46659));
    Odrv12 I__10680 (
            .O(N__46659),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    InMux I__10679 (
            .O(N__46656),
            .I(N__46653));
    LocalMux I__10678 (
            .O(N__46653),
            .I(N__46650));
    Span4Mux_v I__10677 (
            .O(N__46650),
            .I(N__46647));
    Odrv4 I__10676 (
            .O(N__46647),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__10675 (
            .O(N__46644),
            .I(N__46641));
    LocalMux I__10674 (
            .O(N__46641),
            .I(N__46638));
    Span4Mux_h I__10673 (
            .O(N__46638),
            .I(N__46635));
    Odrv4 I__10672 (
            .O(N__46635),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__10671 (
            .O(N__46632),
            .I(N__46627));
    InMux I__10670 (
            .O(N__46631),
            .I(N__46622));
    InMux I__10669 (
            .O(N__46630),
            .I(N__46622));
    LocalMux I__10668 (
            .O(N__46627),
            .I(elapsed_time_ns_1_RNINBNQL1_0_6));
    LocalMux I__10667 (
            .O(N__46622),
            .I(elapsed_time_ns_1_RNINBNQL1_0_6));
    InMux I__10666 (
            .O(N__46617),
            .I(N__46614));
    LocalMux I__10665 (
            .O(N__46614),
            .I(N__46611));
    Span4Mux_h I__10664 (
            .O(N__46611),
            .I(N__46608));
    Odrv4 I__10663 (
            .O(N__46608),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    InMux I__10662 (
            .O(N__46605),
            .I(bfn_18_18_0_));
    InMux I__10661 (
            .O(N__46602),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CascadeMux I__10660 (
            .O(N__46599),
            .I(N__46596));
    InMux I__10659 (
            .O(N__46596),
            .I(N__46591));
    InMux I__10658 (
            .O(N__46595),
            .I(N__46588));
    InMux I__10657 (
            .O(N__46594),
            .I(N__46585));
    LocalMux I__10656 (
            .O(N__46591),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__10655 (
            .O(N__46588),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__10654 (
            .O(N__46585),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__10653 (
            .O(N__46578),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    CascadeMux I__10652 (
            .O(N__46575),
            .I(N__46572));
    InMux I__10651 (
            .O(N__46572),
            .I(N__46567));
    InMux I__10650 (
            .O(N__46571),
            .I(N__46564));
    InMux I__10649 (
            .O(N__46570),
            .I(N__46561));
    LocalMux I__10648 (
            .O(N__46567),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__10647 (
            .O(N__46564),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__10646 (
            .O(N__46561),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__10645 (
            .O(N__46554),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    CascadeMux I__10644 (
            .O(N__46551),
            .I(N__46548));
    InMux I__10643 (
            .O(N__46548),
            .I(N__46544));
    InMux I__10642 (
            .O(N__46547),
            .I(N__46541));
    LocalMux I__10641 (
            .O(N__46544),
            .I(N__46538));
    LocalMux I__10640 (
            .O(N__46541),
            .I(N__46533));
    Span4Mux_v I__10639 (
            .O(N__46538),
            .I(N__46530));
    InMux I__10638 (
            .O(N__46537),
            .I(N__46525));
    InMux I__10637 (
            .O(N__46536),
            .I(N__46525));
    Odrv4 I__10636 (
            .O(N__46533),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    Odrv4 I__10635 (
            .O(N__46530),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    LocalMux I__10634 (
            .O(N__46525),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    InMux I__10633 (
            .O(N__46518),
            .I(N__46515));
    LocalMux I__10632 (
            .O(N__46515),
            .I(N__46512));
    Span4Mux_v I__10631 (
            .O(N__46512),
            .I(N__46509));
    Span4Mux_h I__10630 (
            .O(N__46509),
            .I(N__46506));
    Odrv4 I__10629 (
            .O(N__46506),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    InMux I__10628 (
            .O(N__46503),
            .I(N__46500));
    LocalMux I__10627 (
            .O(N__46500),
            .I(N__46497));
    Span4Mux_v I__10626 (
            .O(N__46497),
            .I(N__46494));
    Span4Mux_h I__10625 (
            .O(N__46494),
            .I(N__46491));
    Span4Mux_h I__10624 (
            .O(N__46491),
            .I(N__46488));
    Odrv4 I__10623 (
            .O(N__46488),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    InMux I__10622 (
            .O(N__46485),
            .I(N__46481));
    InMux I__10621 (
            .O(N__46484),
            .I(N__46477));
    LocalMux I__10620 (
            .O(N__46481),
            .I(N__46474));
    InMux I__10619 (
            .O(N__46480),
            .I(N__46469));
    LocalMux I__10618 (
            .O(N__46477),
            .I(N__46466));
    Span4Mux_v I__10617 (
            .O(N__46474),
            .I(N__46463));
    InMux I__10616 (
            .O(N__46473),
            .I(N__46460));
    InMux I__10615 (
            .O(N__46472),
            .I(N__46457));
    LocalMux I__10614 (
            .O(N__46469),
            .I(elapsed_time_ns_1_RNI8765M1_0_16));
    Odrv12 I__10613 (
            .O(N__46466),
            .I(elapsed_time_ns_1_RNI8765M1_0_16));
    Odrv4 I__10612 (
            .O(N__46463),
            .I(elapsed_time_ns_1_RNI8765M1_0_16));
    LocalMux I__10611 (
            .O(N__46460),
            .I(elapsed_time_ns_1_RNI8765M1_0_16));
    LocalMux I__10610 (
            .O(N__46457),
            .I(elapsed_time_ns_1_RNI8765M1_0_16));
    CascadeMux I__10609 (
            .O(N__46446),
            .I(N__46442));
    InMux I__10608 (
            .O(N__46445),
            .I(N__46437));
    InMux I__10607 (
            .O(N__46442),
            .I(N__46437));
    LocalMux I__10606 (
            .O(N__46437),
            .I(N__46434));
    Span4Mux_h I__10605 (
            .O(N__46434),
            .I(N__46431));
    Odrv4 I__10604 (
            .O(N__46431),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    InMux I__10603 (
            .O(N__46428),
            .I(N__46424));
    InMux I__10602 (
            .O(N__46427),
            .I(N__46419));
    LocalMux I__10601 (
            .O(N__46424),
            .I(N__46416));
    InMux I__10600 (
            .O(N__46423),
            .I(N__46413));
    InMux I__10599 (
            .O(N__46422),
            .I(N__46410));
    LocalMux I__10598 (
            .O(N__46419),
            .I(elapsed_time_ns_1_RNIK8NQL1_0_3));
    Odrv4 I__10597 (
            .O(N__46416),
            .I(elapsed_time_ns_1_RNIK8NQL1_0_3));
    LocalMux I__10596 (
            .O(N__46413),
            .I(elapsed_time_ns_1_RNIK8NQL1_0_3));
    LocalMux I__10595 (
            .O(N__46410),
            .I(elapsed_time_ns_1_RNIK8NQL1_0_3));
    InMux I__10594 (
            .O(N__46401),
            .I(N__46396));
    InMux I__10593 (
            .O(N__46400),
            .I(N__46391));
    InMux I__10592 (
            .O(N__46399),
            .I(N__46391));
    LocalMux I__10591 (
            .O(N__46396),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    LocalMux I__10590 (
            .O(N__46391),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    CascadeMux I__10589 (
            .O(N__46386),
            .I(N__46383));
    InMux I__10588 (
            .O(N__46383),
            .I(N__46379));
    InMux I__10587 (
            .O(N__46382),
            .I(N__46376));
    LocalMux I__10586 (
            .O(N__46379),
            .I(N__46373));
    LocalMux I__10585 (
            .O(N__46376),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ));
    Odrv4 I__10584 (
            .O(N__46373),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ));
    InMux I__10583 (
            .O(N__46368),
            .I(N__46359));
    InMux I__10582 (
            .O(N__46367),
            .I(N__46359));
    InMux I__10581 (
            .O(N__46366),
            .I(N__46359));
    LocalMux I__10580 (
            .O(N__46359),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2 ));
    InMux I__10579 (
            .O(N__46356),
            .I(N__46353));
    LocalMux I__10578 (
            .O(N__46353),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1 ));
    InMux I__10577 (
            .O(N__46350),
            .I(N__46347));
    LocalMux I__10576 (
            .O(N__46347),
            .I(N__46341));
    InMux I__10575 (
            .O(N__46346),
            .I(N__46338));
    InMux I__10574 (
            .O(N__46345),
            .I(N__46333));
    InMux I__10573 (
            .O(N__46344),
            .I(N__46333));
    Odrv4 I__10572 (
            .O(N__46341),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    LocalMux I__10571 (
            .O(N__46338),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    LocalMux I__10570 (
            .O(N__46333),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    CascadeMux I__10569 (
            .O(N__46326),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_ ));
    CascadeMux I__10568 (
            .O(N__46323),
            .I(elapsed_time_ns_1_RNINBNQL1_0_6_cascade_));
    InMux I__10567 (
            .O(N__46320),
            .I(N__46317));
    LocalMux I__10566 (
            .O(N__46317),
            .I(N__46314));
    Span4Mux_v I__10565 (
            .O(N__46314),
            .I(N__46311));
    Span4Mux_h I__10564 (
            .O(N__46311),
            .I(N__46307));
    InMux I__10563 (
            .O(N__46310),
            .I(N__46304));
    Odrv4 I__10562 (
            .O(N__46307),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2 ));
    LocalMux I__10561 (
            .O(N__46304),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2 ));
    CascadeMux I__10560 (
            .O(N__46299),
            .I(N__46295));
    CascadeMux I__10559 (
            .O(N__46298),
            .I(N__46291));
    InMux I__10558 (
            .O(N__46295),
            .I(N__46284));
    InMux I__10557 (
            .O(N__46294),
            .I(N__46284));
    InMux I__10556 (
            .O(N__46291),
            .I(N__46284));
    LocalMux I__10555 (
            .O(N__46284),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ));
    CascadeMux I__10554 (
            .O(N__46281),
            .I(N__46278));
    InMux I__10553 (
            .O(N__46278),
            .I(N__46274));
    CascadeMux I__10552 (
            .O(N__46277),
            .I(N__46270));
    LocalMux I__10551 (
            .O(N__46274),
            .I(N__46266));
    CascadeMux I__10550 (
            .O(N__46273),
            .I(N__46263));
    InMux I__10549 (
            .O(N__46270),
            .I(N__46258));
    InMux I__10548 (
            .O(N__46269),
            .I(N__46258));
    Span4Mux_v I__10547 (
            .O(N__46266),
            .I(N__46255));
    InMux I__10546 (
            .O(N__46263),
            .I(N__46252));
    LocalMux I__10545 (
            .O(N__46258),
            .I(N__46249));
    Span4Mux_h I__10544 (
            .O(N__46255),
            .I(N__46246));
    LocalMux I__10543 (
            .O(N__46252),
            .I(N__46241));
    Span4Mux_v I__10542 (
            .O(N__46249),
            .I(N__46241));
    Odrv4 I__10541 (
            .O(N__46246),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__10540 (
            .O(N__46241),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__10539 (
            .O(N__46236),
            .I(N__46233));
    LocalMux I__10538 (
            .O(N__46233),
            .I(N__46228));
    InMux I__10537 (
            .O(N__46232),
            .I(N__46225));
    InMux I__10536 (
            .O(N__46231),
            .I(N__46222));
    Odrv4 I__10535 (
            .O(N__46228),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__10534 (
            .O(N__46225),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__10533 (
            .O(N__46222),
            .I(\current_shift_inst.un4_control_input1_23 ));
    CascadeMux I__10532 (
            .O(N__46215),
            .I(N__46212));
    InMux I__10531 (
            .O(N__46212),
            .I(N__46209));
    LocalMux I__10530 (
            .O(N__46209),
            .I(N__46206));
    Span4Mux_v I__10529 (
            .O(N__46206),
            .I(N__46203));
    Odrv4 I__10528 (
            .O(N__46203),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__10527 (
            .O(N__46200),
            .I(N__46197));
    LocalMux I__10526 (
            .O(N__46197),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    CascadeMux I__10525 (
            .O(N__46194),
            .I(N__46190));
    InMux I__10524 (
            .O(N__46193),
            .I(N__46186));
    InMux I__10523 (
            .O(N__46190),
            .I(N__46183));
    InMux I__10522 (
            .O(N__46189),
            .I(N__46180));
    LocalMux I__10521 (
            .O(N__46186),
            .I(N__46177));
    LocalMux I__10520 (
            .O(N__46183),
            .I(N__46174));
    LocalMux I__10519 (
            .O(N__46180),
            .I(N__46171));
    Span4Mux_v I__10518 (
            .O(N__46177),
            .I(N__46166));
    Span4Mux_h I__10517 (
            .O(N__46174),
            .I(N__46166));
    Span4Mux_v I__10516 (
            .O(N__46171),
            .I(N__46163));
    Span4Mux_h I__10515 (
            .O(N__46166),
            .I(N__46159));
    Span4Mux_h I__10514 (
            .O(N__46163),
            .I(N__46156));
    InMux I__10513 (
            .O(N__46162),
            .I(N__46153));
    Odrv4 I__10512 (
            .O(N__46159),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__10511 (
            .O(N__46156),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__10510 (
            .O(N__46153),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__10509 (
            .O(N__46146),
            .I(N__46143));
    LocalMux I__10508 (
            .O(N__46143),
            .I(N__46140));
    Span4Mux_v I__10507 (
            .O(N__46140),
            .I(N__46135));
    InMux I__10506 (
            .O(N__46139),
            .I(N__46132));
    InMux I__10505 (
            .O(N__46138),
            .I(N__46129));
    Odrv4 I__10504 (
            .O(N__46135),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__10503 (
            .O(N__46132),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__10502 (
            .O(N__46129),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__10501 (
            .O(N__46122),
            .I(N__46119));
    LocalMux I__10500 (
            .O(N__46119),
            .I(N__46116));
    Odrv4 I__10499 (
            .O(N__46116),
            .I(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ));
    CascadeMux I__10498 (
            .O(N__46113),
            .I(N__46109));
    CascadeMux I__10497 (
            .O(N__46112),
            .I(N__46106));
    InMux I__10496 (
            .O(N__46109),
            .I(N__46102));
    InMux I__10495 (
            .O(N__46106),
            .I(N__46099));
    InMux I__10494 (
            .O(N__46105),
            .I(N__46096));
    LocalMux I__10493 (
            .O(N__46102),
            .I(N__46092));
    LocalMux I__10492 (
            .O(N__46099),
            .I(N__46089));
    LocalMux I__10491 (
            .O(N__46096),
            .I(N__46086));
    InMux I__10490 (
            .O(N__46095),
            .I(N__46083));
    Span4Mux_h I__10489 (
            .O(N__46092),
            .I(N__46080));
    Span4Mux_v I__10488 (
            .O(N__46089),
            .I(N__46077));
    Span4Mux_h I__10487 (
            .O(N__46086),
            .I(N__46074));
    LocalMux I__10486 (
            .O(N__46083),
            .I(N__46071));
    Span4Mux_h I__10485 (
            .O(N__46080),
            .I(N__46068));
    Span4Mux_h I__10484 (
            .O(N__46077),
            .I(N__46063));
    Span4Mux_h I__10483 (
            .O(N__46074),
            .I(N__46063));
    Odrv12 I__10482 (
            .O(N__46071),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__10481 (
            .O(N__46068),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__10480 (
            .O(N__46063),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__10479 (
            .O(N__46056),
            .I(N__46053));
    LocalMux I__10478 (
            .O(N__46053),
            .I(N__46049));
    InMux I__10477 (
            .O(N__46052),
            .I(N__46046));
    Span4Mux_v I__10476 (
            .O(N__46049),
            .I(N__46042));
    LocalMux I__10475 (
            .O(N__46046),
            .I(N__46039));
    InMux I__10474 (
            .O(N__46045),
            .I(N__46036));
    Odrv4 I__10473 (
            .O(N__46042),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__10472 (
            .O(N__46039),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__10471 (
            .O(N__46036),
            .I(\current_shift_inst.un4_control_input1_15 ));
    CascadeMux I__10470 (
            .O(N__46029),
            .I(N__46026));
    InMux I__10469 (
            .O(N__46026),
            .I(N__46023));
    LocalMux I__10468 (
            .O(N__46023),
            .I(N__46020));
    Span4Mux_h I__10467 (
            .O(N__46020),
            .I(N__46017));
    Odrv4 I__10466 (
            .O(N__46017),
            .I(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ));
    CascadeMux I__10465 (
            .O(N__46014),
            .I(N__45989));
    CascadeMux I__10464 (
            .O(N__46013),
            .I(N__45983));
    CascadeMux I__10463 (
            .O(N__46012),
            .I(N__45977));
    InMux I__10462 (
            .O(N__46011),
            .I(N__45965));
    InMux I__10461 (
            .O(N__46010),
            .I(N__45965));
    InMux I__10460 (
            .O(N__46009),
            .I(N__45965));
    InMux I__10459 (
            .O(N__46008),
            .I(N__45965));
    InMux I__10458 (
            .O(N__46007),
            .I(N__45956));
    InMux I__10457 (
            .O(N__46006),
            .I(N__45956));
    InMux I__10456 (
            .O(N__46005),
            .I(N__45956));
    InMux I__10455 (
            .O(N__46004),
            .I(N__45956));
    CascadeMux I__10454 (
            .O(N__46003),
            .I(N__45949));
    CascadeMux I__10453 (
            .O(N__46002),
            .I(N__45936));
    CascadeMux I__10452 (
            .O(N__46001),
            .I(N__45932));
    CascadeMux I__10451 (
            .O(N__46000),
            .I(N__45928));
    CascadeMux I__10450 (
            .O(N__45999),
            .I(N__45924));
    CascadeMux I__10449 (
            .O(N__45998),
            .I(N__45920));
    CascadeMux I__10448 (
            .O(N__45997),
            .I(N__45916));
    CascadeMux I__10447 (
            .O(N__45996),
            .I(N__45912));
    CascadeMux I__10446 (
            .O(N__45995),
            .I(N__45897));
    CascadeMux I__10445 (
            .O(N__45994),
            .I(N__45893));
    CascadeMux I__10444 (
            .O(N__45993),
            .I(N__45889));
    InMux I__10443 (
            .O(N__45992),
            .I(N__45877));
    InMux I__10442 (
            .O(N__45989),
            .I(N__45877));
    InMux I__10441 (
            .O(N__45988),
            .I(N__45871));
    InMux I__10440 (
            .O(N__45987),
            .I(N__45864));
    InMux I__10439 (
            .O(N__45986),
            .I(N__45864));
    InMux I__10438 (
            .O(N__45983),
            .I(N__45864));
    InMux I__10437 (
            .O(N__45982),
            .I(N__45853));
    InMux I__10436 (
            .O(N__45981),
            .I(N__45853));
    InMux I__10435 (
            .O(N__45980),
            .I(N__45853));
    InMux I__10434 (
            .O(N__45977),
            .I(N__45853));
    InMux I__10433 (
            .O(N__45976),
            .I(N__45853));
    CascadeMux I__10432 (
            .O(N__45975),
            .I(N__45849));
    CascadeMux I__10431 (
            .O(N__45974),
            .I(N__45845));
    LocalMux I__10430 (
            .O(N__45965),
            .I(N__45835));
    LocalMux I__10429 (
            .O(N__45956),
            .I(N__45835));
    InMux I__10428 (
            .O(N__45955),
            .I(N__45822));
    InMux I__10427 (
            .O(N__45954),
            .I(N__45822));
    InMux I__10426 (
            .O(N__45953),
            .I(N__45822));
    InMux I__10425 (
            .O(N__45952),
            .I(N__45822));
    InMux I__10424 (
            .O(N__45949),
            .I(N__45822));
    InMux I__10423 (
            .O(N__45948),
            .I(N__45822));
    InMux I__10422 (
            .O(N__45947),
            .I(N__45811));
    InMux I__10421 (
            .O(N__45946),
            .I(N__45811));
    InMux I__10420 (
            .O(N__45945),
            .I(N__45811));
    InMux I__10419 (
            .O(N__45944),
            .I(N__45811));
    InMux I__10418 (
            .O(N__45943),
            .I(N__45811));
    InMux I__10417 (
            .O(N__45942),
            .I(N__45806));
    InMux I__10416 (
            .O(N__45941),
            .I(N__45806));
    InMux I__10415 (
            .O(N__45940),
            .I(N__45784));
    InMux I__10414 (
            .O(N__45939),
            .I(N__45784));
    InMux I__10413 (
            .O(N__45936),
            .I(N__45784));
    InMux I__10412 (
            .O(N__45935),
            .I(N__45784));
    InMux I__10411 (
            .O(N__45932),
            .I(N__45784));
    InMux I__10410 (
            .O(N__45931),
            .I(N__45784));
    InMux I__10409 (
            .O(N__45928),
            .I(N__45784));
    InMux I__10408 (
            .O(N__45927),
            .I(N__45784));
    InMux I__10407 (
            .O(N__45924),
            .I(N__45767));
    InMux I__10406 (
            .O(N__45923),
            .I(N__45767));
    InMux I__10405 (
            .O(N__45920),
            .I(N__45767));
    InMux I__10404 (
            .O(N__45919),
            .I(N__45767));
    InMux I__10403 (
            .O(N__45916),
            .I(N__45767));
    InMux I__10402 (
            .O(N__45915),
            .I(N__45767));
    InMux I__10401 (
            .O(N__45912),
            .I(N__45767));
    InMux I__10400 (
            .O(N__45911),
            .I(N__45767));
    CascadeMux I__10399 (
            .O(N__45910),
            .I(N__45764));
    CascadeMux I__10398 (
            .O(N__45909),
            .I(N__45760));
    CascadeMux I__10397 (
            .O(N__45908),
            .I(N__45756));
    CascadeMux I__10396 (
            .O(N__45907),
            .I(N__45752));
    CascadeMux I__10395 (
            .O(N__45906),
            .I(N__45744));
    CascadeMux I__10394 (
            .O(N__45905),
            .I(N__45740));
    CascadeMux I__10393 (
            .O(N__45904),
            .I(N__45736));
    CascadeMux I__10392 (
            .O(N__45903),
            .I(N__45732));
    CascadeMux I__10391 (
            .O(N__45902),
            .I(N__45728));
    CascadeMux I__10390 (
            .O(N__45901),
            .I(N__45724));
    CascadeMux I__10389 (
            .O(N__45900),
            .I(N__45720));
    InMux I__10388 (
            .O(N__45897),
            .I(N__45706));
    InMux I__10387 (
            .O(N__45896),
            .I(N__45706));
    InMux I__10386 (
            .O(N__45893),
            .I(N__45706));
    InMux I__10385 (
            .O(N__45892),
            .I(N__45706));
    InMux I__10384 (
            .O(N__45889),
            .I(N__45706));
    InMux I__10383 (
            .O(N__45888),
            .I(N__45706));
    InMux I__10382 (
            .O(N__45887),
            .I(N__45697));
    InMux I__10381 (
            .O(N__45886),
            .I(N__45697));
    InMux I__10380 (
            .O(N__45885),
            .I(N__45697));
    InMux I__10379 (
            .O(N__45884),
            .I(N__45697));
    InMux I__10378 (
            .O(N__45883),
            .I(N__45692));
    InMux I__10377 (
            .O(N__45882),
            .I(N__45692));
    LocalMux I__10376 (
            .O(N__45877),
            .I(N__45689));
    InMux I__10375 (
            .O(N__45876),
            .I(N__45686));
    CascadeMux I__10374 (
            .O(N__45875),
            .I(N__45682));
    CascadeMux I__10373 (
            .O(N__45874),
            .I(N__45676));
    LocalMux I__10372 (
            .O(N__45871),
            .I(N__45667));
    LocalMux I__10371 (
            .O(N__45864),
            .I(N__45667));
    LocalMux I__10370 (
            .O(N__45853),
            .I(N__45664));
    InMux I__10369 (
            .O(N__45852),
            .I(N__45653));
    InMux I__10368 (
            .O(N__45849),
            .I(N__45653));
    InMux I__10367 (
            .O(N__45848),
            .I(N__45653));
    InMux I__10366 (
            .O(N__45845),
            .I(N__45653));
    InMux I__10365 (
            .O(N__45844),
            .I(N__45653));
    CascadeMux I__10364 (
            .O(N__45843),
            .I(N__45650));
    CascadeMux I__10363 (
            .O(N__45842),
            .I(N__45646));
    CascadeMux I__10362 (
            .O(N__45841),
            .I(N__45642));
    CascadeMux I__10361 (
            .O(N__45840),
            .I(N__45638));
    Span4Mux_v I__10360 (
            .O(N__45835),
            .I(N__45628));
    LocalMux I__10359 (
            .O(N__45822),
            .I(N__45628));
    LocalMux I__10358 (
            .O(N__45811),
            .I(N__45628));
    LocalMux I__10357 (
            .O(N__45806),
            .I(N__45628));
    InMux I__10356 (
            .O(N__45805),
            .I(N__45617));
    InMux I__10355 (
            .O(N__45804),
            .I(N__45617));
    InMux I__10354 (
            .O(N__45803),
            .I(N__45617));
    InMux I__10353 (
            .O(N__45802),
            .I(N__45617));
    InMux I__10352 (
            .O(N__45801),
            .I(N__45617));
    LocalMux I__10351 (
            .O(N__45784),
            .I(N__45612));
    LocalMux I__10350 (
            .O(N__45767),
            .I(N__45612));
    InMux I__10349 (
            .O(N__45764),
            .I(N__45595));
    InMux I__10348 (
            .O(N__45763),
            .I(N__45595));
    InMux I__10347 (
            .O(N__45760),
            .I(N__45595));
    InMux I__10346 (
            .O(N__45759),
            .I(N__45595));
    InMux I__10345 (
            .O(N__45756),
            .I(N__45595));
    InMux I__10344 (
            .O(N__45755),
            .I(N__45595));
    InMux I__10343 (
            .O(N__45752),
            .I(N__45595));
    InMux I__10342 (
            .O(N__45751),
            .I(N__45595));
    CascadeMux I__10341 (
            .O(N__45750),
            .I(N__45592));
    CascadeMux I__10340 (
            .O(N__45749),
            .I(N__45588));
    CascadeMux I__10339 (
            .O(N__45748),
            .I(N__45584));
    InMux I__10338 (
            .O(N__45747),
            .I(N__45568));
    InMux I__10337 (
            .O(N__45744),
            .I(N__45568));
    InMux I__10336 (
            .O(N__45743),
            .I(N__45568));
    InMux I__10335 (
            .O(N__45740),
            .I(N__45568));
    InMux I__10334 (
            .O(N__45739),
            .I(N__45568));
    InMux I__10333 (
            .O(N__45736),
            .I(N__45568));
    InMux I__10332 (
            .O(N__45735),
            .I(N__45568));
    InMux I__10331 (
            .O(N__45732),
            .I(N__45551));
    InMux I__10330 (
            .O(N__45731),
            .I(N__45551));
    InMux I__10329 (
            .O(N__45728),
            .I(N__45551));
    InMux I__10328 (
            .O(N__45727),
            .I(N__45551));
    InMux I__10327 (
            .O(N__45724),
            .I(N__45551));
    InMux I__10326 (
            .O(N__45723),
            .I(N__45551));
    InMux I__10325 (
            .O(N__45720),
            .I(N__45551));
    InMux I__10324 (
            .O(N__45719),
            .I(N__45551));
    LocalMux I__10323 (
            .O(N__45706),
            .I(N__45548));
    LocalMux I__10322 (
            .O(N__45697),
            .I(N__45543));
    LocalMux I__10321 (
            .O(N__45692),
            .I(N__45543));
    Span4Mux_h I__10320 (
            .O(N__45689),
            .I(N__45538));
    LocalMux I__10319 (
            .O(N__45686),
            .I(N__45538));
    InMux I__10318 (
            .O(N__45685),
            .I(N__45523));
    InMux I__10317 (
            .O(N__45682),
            .I(N__45523));
    InMux I__10316 (
            .O(N__45681),
            .I(N__45523));
    InMux I__10315 (
            .O(N__45680),
            .I(N__45523));
    InMux I__10314 (
            .O(N__45679),
            .I(N__45523));
    InMux I__10313 (
            .O(N__45676),
            .I(N__45523));
    InMux I__10312 (
            .O(N__45675),
            .I(N__45523));
    InMux I__10311 (
            .O(N__45674),
            .I(N__45516));
    InMux I__10310 (
            .O(N__45673),
            .I(N__45516));
    InMux I__10309 (
            .O(N__45672),
            .I(N__45516));
    Span4Mux_v I__10308 (
            .O(N__45667),
            .I(N__45509));
    Span4Mux_v I__10307 (
            .O(N__45664),
            .I(N__45509));
    LocalMux I__10306 (
            .O(N__45653),
            .I(N__45509));
    InMux I__10305 (
            .O(N__45650),
            .I(N__45492));
    InMux I__10304 (
            .O(N__45649),
            .I(N__45492));
    InMux I__10303 (
            .O(N__45646),
            .I(N__45492));
    InMux I__10302 (
            .O(N__45645),
            .I(N__45492));
    InMux I__10301 (
            .O(N__45642),
            .I(N__45492));
    InMux I__10300 (
            .O(N__45641),
            .I(N__45492));
    InMux I__10299 (
            .O(N__45638),
            .I(N__45492));
    InMux I__10298 (
            .O(N__45637),
            .I(N__45492));
    Span4Mux_v I__10297 (
            .O(N__45628),
            .I(N__45483));
    LocalMux I__10296 (
            .O(N__45617),
            .I(N__45483));
    Span4Mux_v I__10295 (
            .O(N__45612),
            .I(N__45483));
    LocalMux I__10294 (
            .O(N__45595),
            .I(N__45483));
    InMux I__10293 (
            .O(N__45592),
            .I(N__45470));
    InMux I__10292 (
            .O(N__45591),
            .I(N__45470));
    InMux I__10291 (
            .O(N__45588),
            .I(N__45470));
    InMux I__10290 (
            .O(N__45587),
            .I(N__45470));
    InMux I__10289 (
            .O(N__45584),
            .I(N__45470));
    InMux I__10288 (
            .O(N__45583),
            .I(N__45470));
    LocalMux I__10287 (
            .O(N__45568),
            .I(N__45463));
    LocalMux I__10286 (
            .O(N__45551),
            .I(N__45463));
    Span4Mux_h I__10285 (
            .O(N__45548),
            .I(N__45463));
    Odrv12 I__10284 (
            .O(N__45543),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10283 (
            .O(N__45538),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10282 (
            .O(N__45523),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10281 (
            .O(N__45516),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10280 (
            .O(N__45509),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10279 (
            .O(N__45492),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10278 (
            .O(N__45483),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10277 (
            .O(N__45470),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10276 (
            .O(N__45463),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__10275 (
            .O(N__45444),
            .I(N__45400));
    InMux I__10274 (
            .O(N__45443),
            .I(N__45389));
    InMux I__10273 (
            .O(N__45442),
            .I(N__45378));
    InMux I__10272 (
            .O(N__45441),
            .I(N__45378));
    InMux I__10271 (
            .O(N__45440),
            .I(N__45378));
    InMux I__10270 (
            .O(N__45439),
            .I(N__45378));
    InMux I__10269 (
            .O(N__45438),
            .I(N__45378));
    InMux I__10268 (
            .O(N__45437),
            .I(N__45365));
    InMux I__10267 (
            .O(N__45436),
            .I(N__45365));
    InMux I__10266 (
            .O(N__45435),
            .I(N__45365));
    InMux I__10265 (
            .O(N__45434),
            .I(N__45365));
    InMux I__10264 (
            .O(N__45433),
            .I(N__45365));
    InMux I__10263 (
            .O(N__45432),
            .I(N__45365));
    InMux I__10262 (
            .O(N__45431),
            .I(N__45355));
    InMux I__10261 (
            .O(N__45430),
            .I(N__45355));
    InMux I__10260 (
            .O(N__45429),
            .I(N__45355));
    InMux I__10259 (
            .O(N__45428),
            .I(N__45355));
    InMux I__10258 (
            .O(N__45427),
            .I(N__45346));
    InMux I__10257 (
            .O(N__45426),
            .I(N__45346));
    InMux I__10256 (
            .O(N__45425),
            .I(N__45346));
    InMux I__10255 (
            .O(N__45424),
            .I(N__45346));
    InMux I__10254 (
            .O(N__45423),
            .I(N__45333));
    InMux I__10253 (
            .O(N__45422),
            .I(N__45333));
    InMux I__10252 (
            .O(N__45421),
            .I(N__45324));
    InMux I__10251 (
            .O(N__45420),
            .I(N__45324));
    InMux I__10250 (
            .O(N__45419),
            .I(N__45324));
    InMux I__10249 (
            .O(N__45418),
            .I(N__45324));
    InMux I__10248 (
            .O(N__45417),
            .I(N__45313));
    InMux I__10247 (
            .O(N__45416),
            .I(N__45313));
    InMux I__10246 (
            .O(N__45415),
            .I(N__45313));
    InMux I__10245 (
            .O(N__45414),
            .I(N__45313));
    InMux I__10244 (
            .O(N__45413),
            .I(N__45313));
    InMux I__10243 (
            .O(N__45412),
            .I(N__45306));
    InMux I__10242 (
            .O(N__45411),
            .I(N__45306));
    InMux I__10241 (
            .O(N__45410),
            .I(N__45306));
    InMux I__10240 (
            .O(N__45409),
            .I(N__45303));
    InMux I__10239 (
            .O(N__45408),
            .I(N__45286));
    InMux I__10238 (
            .O(N__45407),
            .I(N__45286));
    InMux I__10237 (
            .O(N__45406),
            .I(N__45286));
    InMux I__10236 (
            .O(N__45405),
            .I(N__45286));
    InMux I__10235 (
            .O(N__45404),
            .I(N__45286));
    InMux I__10234 (
            .O(N__45403),
            .I(N__45283));
    InMux I__10233 (
            .O(N__45400),
            .I(N__45268));
    InMux I__10232 (
            .O(N__45399),
            .I(N__45268));
    InMux I__10231 (
            .O(N__45398),
            .I(N__45268));
    InMux I__10230 (
            .O(N__45397),
            .I(N__45268));
    InMux I__10229 (
            .O(N__45396),
            .I(N__45268));
    InMux I__10228 (
            .O(N__45395),
            .I(N__45268));
    InMux I__10227 (
            .O(N__45394),
            .I(N__45268));
    InMux I__10226 (
            .O(N__45393),
            .I(N__45263));
    InMux I__10225 (
            .O(N__45392),
            .I(N__45260));
    LocalMux I__10224 (
            .O(N__45389),
            .I(N__45257));
    LocalMux I__10223 (
            .O(N__45378),
            .I(N__45252));
    LocalMux I__10222 (
            .O(N__45365),
            .I(N__45252));
    CascadeMux I__10221 (
            .O(N__45364),
            .I(N__45246));
    LocalMux I__10220 (
            .O(N__45355),
            .I(N__45242));
    LocalMux I__10219 (
            .O(N__45346),
            .I(N__45239));
    InMux I__10218 (
            .O(N__45345),
            .I(N__45236));
    InMux I__10217 (
            .O(N__45344),
            .I(N__45221));
    InMux I__10216 (
            .O(N__45343),
            .I(N__45221));
    InMux I__10215 (
            .O(N__45342),
            .I(N__45221));
    InMux I__10214 (
            .O(N__45341),
            .I(N__45221));
    InMux I__10213 (
            .O(N__45340),
            .I(N__45221));
    InMux I__10212 (
            .O(N__45339),
            .I(N__45221));
    InMux I__10211 (
            .O(N__45338),
            .I(N__45221));
    LocalMux I__10210 (
            .O(N__45333),
            .I(N__45216));
    LocalMux I__10209 (
            .O(N__45324),
            .I(N__45216));
    LocalMux I__10208 (
            .O(N__45313),
            .I(N__45213));
    LocalMux I__10207 (
            .O(N__45306),
            .I(N__45208));
    LocalMux I__10206 (
            .O(N__45303),
            .I(N__45208));
    InMux I__10205 (
            .O(N__45302),
            .I(N__45195));
    InMux I__10204 (
            .O(N__45301),
            .I(N__45195));
    InMux I__10203 (
            .O(N__45300),
            .I(N__45195));
    InMux I__10202 (
            .O(N__45299),
            .I(N__45195));
    InMux I__10201 (
            .O(N__45298),
            .I(N__45195));
    InMux I__10200 (
            .O(N__45297),
            .I(N__45195));
    LocalMux I__10199 (
            .O(N__45286),
            .I(N__45192));
    LocalMux I__10198 (
            .O(N__45283),
            .I(N__45187));
    LocalMux I__10197 (
            .O(N__45268),
            .I(N__45187));
    InMux I__10196 (
            .O(N__45267),
            .I(N__45182));
    InMux I__10195 (
            .O(N__45266),
            .I(N__45182));
    LocalMux I__10194 (
            .O(N__45263),
            .I(N__45173));
    LocalMux I__10193 (
            .O(N__45260),
            .I(N__45173));
    Span4Mux_v I__10192 (
            .O(N__45257),
            .I(N__45173));
    Span4Mux_v I__10191 (
            .O(N__45252),
            .I(N__45173));
    InMux I__10190 (
            .O(N__45251),
            .I(N__45162));
    InMux I__10189 (
            .O(N__45250),
            .I(N__45162));
    InMux I__10188 (
            .O(N__45249),
            .I(N__45162));
    InMux I__10187 (
            .O(N__45246),
            .I(N__45162));
    InMux I__10186 (
            .O(N__45245),
            .I(N__45162));
    Span4Mux_h I__10185 (
            .O(N__45242),
            .I(N__45159));
    Span4Mux_v I__10184 (
            .O(N__45239),
            .I(N__45156));
    LocalMux I__10183 (
            .O(N__45236),
            .I(N__45145));
    LocalMux I__10182 (
            .O(N__45221),
            .I(N__45145));
    Span4Mux_v I__10181 (
            .O(N__45216),
            .I(N__45145));
    Span4Mux_h I__10180 (
            .O(N__45213),
            .I(N__45145));
    Span4Mux_v I__10179 (
            .O(N__45208),
            .I(N__45145));
    LocalMux I__10178 (
            .O(N__45195),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10177 (
            .O(N__45192),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10176 (
            .O(N__45187),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10175 (
            .O(N__45182),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10174 (
            .O(N__45173),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10173 (
            .O(N__45162),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10172 (
            .O(N__45159),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10171 (
            .O(N__45156),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10170 (
            .O(N__45145),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__10169 (
            .O(N__45126),
            .I(N__45123));
    InMux I__10168 (
            .O(N__45123),
            .I(N__45119));
    CascadeMux I__10167 (
            .O(N__45122),
            .I(N__45116));
    LocalMux I__10166 (
            .O(N__45119),
            .I(N__45112));
    InMux I__10165 (
            .O(N__45116),
            .I(N__45107));
    InMux I__10164 (
            .O(N__45115),
            .I(N__45107));
    Odrv4 I__10163 (
            .O(N__45112),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__10162 (
            .O(N__45107),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__10161 (
            .O(N__45102),
            .I(N__45096));
    InMux I__10160 (
            .O(N__45101),
            .I(N__45096));
    LocalMux I__10159 (
            .O(N__45096),
            .I(N__45091));
    InMux I__10158 (
            .O(N__45095),
            .I(N__45086));
    InMux I__10157 (
            .O(N__45094),
            .I(N__45086));
    Span4Mux_h I__10156 (
            .O(N__45091),
            .I(N__45083));
    LocalMux I__10155 (
            .O(N__45086),
            .I(N__45080));
    Span4Mux_h I__10154 (
            .O(N__45083),
            .I(N__45077));
    Odrv4 I__10153 (
            .O(N__45080),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__10152 (
            .O(N__45077),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    CascadeMux I__10151 (
            .O(N__45072),
            .I(N__45069));
    InMux I__10150 (
            .O(N__45069),
            .I(N__45066));
    LocalMux I__10149 (
            .O(N__45066),
            .I(N__45063));
    Span4Mux_h I__10148 (
            .O(N__45063),
            .I(N__45060));
    Odrv4 I__10147 (
            .O(N__45060),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__10146 (
            .O(N__45057),
            .I(N__45054));
    LocalMux I__10145 (
            .O(N__45054),
            .I(N__45051));
    Span4Mux_h I__10144 (
            .O(N__45051),
            .I(N__45048));
    Span4Mux_v I__10143 (
            .O(N__45048),
            .I(N__45045));
    Odrv4 I__10142 (
            .O(N__45045),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__10141 (
            .O(N__45042),
            .I(N__45039));
    InMux I__10140 (
            .O(N__45039),
            .I(N__45036));
    LocalMux I__10139 (
            .O(N__45036),
            .I(N__45033));
    Span4Mux_v I__10138 (
            .O(N__45033),
            .I(N__45029));
    InMux I__10137 (
            .O(N__45032),
            .I(N__45026));
    Odrv4 I__10136 (
            .O(N__45029),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    LocalMux I__10135 (
            .O(N__45026),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__10134 (
            .O(N__45021),
            .I(N__45018));
    LocalMux I__10133 (
            .O(N__45018),
            .I(N__45015));
    Span4Mux_h I__10132 (
            .O(N__45015),
            .I(N__45012));
    Span4Mux_h I__10131 (
            .O(N__45012),
            .I(N__45009));
    Odrv4 I__10130 (
            .O(N__45009),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__10129 (
            .O(N__45006),
            .I(N__45003));
    InMux I__10128 (
            .O(N__45003),
            .I(N__44999));
    CascadeMux I__10127 (
            .O(N__45002),
            .I(N__44995));
    LocalMux I__10126 (
            .O(N__44999),
            .I(N__44991));
    InMux I__10125 (
            .O(N__44998),
            .I(N__44988));
    InMux I__10124 (
            .O(N__44995),
            .I(N__44985));
    InMux I__10123 (
            .O(N__44994),
            .I(N__44982));
    Span4Mux_v I__10122 (
            .O(N__44991),
            .I(N__44977));
    LocalMux I__10121 (
            .O(N__44988),
            .I(N__44977));
    LocalMux I__10120 (
            .O(N__44985),
            .I(N__44974));
    LocalMux I__10119 (
            .O(N__44982),
            .I(N__44969));
    Span4Mux_v I__10118 (
            .O(N__44977),
            .I(N__44969));
    Odrv12 I__10117 (
            .O(N__44974),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__10116 (
            .O(N__44969),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__10115 (
            .O(N__44964),
            .I(N__44961));
    LocalMux I__10114 (
            .O(N__44961),
            .I(N__44958));
    Span4Mux_v I__10113 (
            .O(N__44958),
            .I(N__44953));
    InMux I__10112 (
            .O(N__44957),
            .I(N__44950));
    InMux I__10111 (
            .O(N__44956),
            .I(N__44947));
    Odrv4 I__10110 (
            .O(N__44953),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__10109 (
            .O(N__44950),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__10108 (
            .O(N__44947),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__10107 (
            .O(N__44940),
            .I(N__44937));
    LocalMux I__10106 (
            .O(N__44937),
            .I(N__44934));
    Span4Mux_v I__10105 (
            .O(N__44934),
            .I(N__44931));
    Odrv4 I__10104 (
            .O(N__44931),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__10103 (
            .O(N__44928),
            .I(N__44925));
    LocalMux I__10102 (
            .O(N__44925),
            .I(N__44921));
    InMux I__10101 (
            .O(N__44924),
            .I(N__44918));
    Sp12to4 I__10100 (
            .O(N__44921),
            .I(N__44912));
    LocalMux I__10099 (
            .O(N__44918),
            .I(N__44912));
    InMux I__10098 (
            .O(N__44917),
            .I(N__44909));
    Span12Mux_v I__10097 (
            .O(N__44912),
            .I(N__44906));
    LocalMux I__10096 (
            .O(N__44909),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    Odrv12 I__10095 (
            .O(N__44906),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    InMux I__10094 (
            .O(N__44901),
            .I(N__44893));
    InMux I__10093 (
            .O(N__44900),
            .I(N__44893));
    InMux I__10092 (
            .O(N__44899),
            .I(N__44890));
    InMux I__10091 (
            .O(N__44898),
            .I(N__44887));
    LocalMux I__10090 (
            .O(N__44893),
            .I(N__44884));
    LocalMux I__10089 (
            .O(N__44890),
            .I(N__44881));
    LocalMux I__10088 (
            .O(N__44887),
            .I(N__44878));
    Span4Mux_v I__10087 (
            .O(N__44884),
            .I(N__44875));
    Span12Mux_s9_v I__10086 (
            .O(N__44881),
            .I(N__44872));
    Span4Mux_h I__10085 (
            .O(N__44878),
            .I(N__44869));
    Odrv4 I__10084 (
            .O(N__44875),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv12 I__10083 (
            .O(N__44872),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv4 I__10082 (
            .O(N__44869),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    CascadeMux I__10081 (
            .O(N__44862),
            .I(N__44859));
    InMux I__10080 (
            .O(N__44859),
            .I(N__44852));
    InMux I__10079 (
            .O(N__44858),
            .I(N__44852));
    InMux I__10078 (
            .O(N__44857),
            .I(N__44849));
    LocalMux I__10077 (
            .O(N__44852),
            .I(N__44846));
    LocalMux I__10076 (
            .O(N__44849),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__10075 (
            .O(N__44846),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__10074 (
            .O(N__44841),
            .I(N__44838));
    LocalMux I__10073 (
            .O(N__44838),
            .I(N__44835));
    Span4Mux_v I__10072 (
            .O(N__44835),
            .I(N__44832));
    Odrv4 I__10071 (
            .O(N__44832),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    CascadeMux I__10070 (
            .O(N__44829),
            .I(N__44826));
    InMux I__10069 (
            .O(N__44826),
            .I(N__44822));
    CascadeMux I__10068 (
            .O(N__44825),
            .I(N__44819));
    LocalMux I__10067 (
            .O(N__44822),
            .I(N__44816));
    InMux I__10066 (
            .O(N__44819),
            .I(N__44813));
    Span4Mux_h I__10065 (
            .O(N__44816),
            .I(N__44809));
    LocalMux I__10064 (
            .O(N__44813),
            .I(N__44806));
    CascadeMux I__10063 (
            .O(N__44812),
            .I(N__44803));
    Span4Mux_v I__10062 (
            .O(N__44809),
            .I(N__44797));
    Span4Mux_h I__10061 (
            .O(N__44806),
            .I(N__44797));
    InMux I__10060 (
            .O(N__44803),
            .I(N__44792));
    InMux I__10059 (
            .O(N__44802),
            .I(N__44792));
    Span4Mux_h I__10058 (
            .O(N__44797),
            .I(N__44789));
    LocalMux I__10057 (
            .O(N__44792),
            .I(N__44786));
    Odrv4 I__10056 (
            .O(N__44789),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__10055 (
            .O(N__44786),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__10054 (
            .O(N__44781),
            .I(N__44778));
    LocalMux I__10053 (
            .O(N__44778),
            .I(N__44775));
    Span4Mux_v I__10052 (
            .O(N__44775),
            .I(N__44770));
    InMux I__10051 (
            .O(N__44774),
            .I(N__44767));
    InMux I__10050 (
            .O(N__44773),
            .I(N__44764));
    Odrv4 I__10049 (
            .O(N__44770),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__10048 (
            .O(N__44767),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__10047 (
            .O(N__44764),
            .I(\current_shift_inst.un4_control_input1_11 ));
    CascadeMux I__10046 (
            .O(N__44757),
            .I(N__44754));
    InMux I__10045 (
            .O(N__44754),
            .I(N__44751));
    LocalMux I__10044 (
            .O(N__44751),
            .I(N__44748));
    Odrv4 I__10043 (
            .O(N__44748),
            .I(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ));
    InMux I__10042 (
            .O(N__44745),
            .I(N__44742));
    LocalMux I__10041 (
            .O(N__44742),
            .I(N__44737));
    InMux I__10040 (
            .O(N__44741),
            .I(N__44734));
    InMux I__10039 (
            .O(N__44740),
            .I(N__44729));
    Span4Mux_v I__10038 (
            .O(N__44737),
            .I(N__44726));
    LocalMux I__10037 (
            .O(N__44734),
            .I(N__44723));
    InMux I__10036 (
            .O(N__44733),
            .I(N__44718));
    InMux I__10035 (
            .O(N__44732),
            .I(N__44718));
    LocalMux I__10034 (
            .O(N__44729),
            .I(N__44715));
    Span4Mux_h I__10033 (
            .O(N__44726),
            .I(N__44712));
    Span4Mux_h I__10032 (
            .O(N__44723),
            .I(N__44709));
    LocalMux I__10031 (
            .O(N__44718),
            .I(N__44706));
    Span4Mux_v I__10030 (
            .O(N__44715),
            .I(N__44701));
    Span4Mux_h I__10029 (
            .O(N__44712),
            .I(N__44701));
    Odrv4 I__10028 (
            .O(N__44709),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__10027 (
            .O(N__44706),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__10026 (
            .O(N__44701),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__10025 (
            .O(N__44694),
            .I(N__44691));
    LocalMux I__10024 (
            .O(N__44691),
            .I(N__44688));
    Span4Mux_h I__10023 (
            .O(N__44688),
            .I(N__44685));
    Span4Mux_h I__10022 (
            .O(N__44685),
            .I(N__44682));
    Span4Mux_h I__10021 (
            .O(N__44682),
            .I(N__44679));
    Odrv4 I__10020 (
            .O(N__44679),
            .I(\current_shift_inst.PI_CTRL.integrator_i_25 ));
    CascadeMux I__10019 (
            .O(N__44676),
            .I(N__44672));
    CascadeMux I__10018 (
            .O(N__44675),
            .I(N__44668));
    InMux I__10017 (
            .O(N__44672),
            .I(N__44665));
    InMux I__10016 (
            .O(N__44671),
            .I(N__44662));
    InMux I__10015 (
            .O(N__44668),
            .I(N__44659));
    LocalMux I__10014 (
            .O(N__44665),
            .I(N__44656));
    LocalMux I__10013 (
            .O(N__44662),
            .I(N__44653));
    LocalMux I__10012 (
            .O(N__44659),
            .I(N__44649));
    Span4Mux_v I__10011 (
            .O(N__44656),
            .I(N__44644));
    Span4Mux_h I__10010 (
            .O(N__44653),
            .I(N__44644));
    InMux I__10009 (
            .O(N__44652),
            .I(N__44641));
    Odrv12 I__10008 (
            .O(N__44649),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__10007 (
            .O(N__44644),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__10006 (
            .O(N__44641),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__10005 (
            .O(N__44634),
            .I(N__44631));
    LocalMux I__10004 (
            .O(N__44631),
            .I(N__44628));
    Span4Mux_h I__10003 (
            .O(N__44628),
            .I(N__44623));
    InMux I__10002 (
            .O(N__44627),
            .I(N__44620));
    InMux I__10001 (
            .O(N__44626),
            .I(N__44617));
    Odrv4 I__10000 (
            .O(N__44623),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__9999 (
            .O(N__44620),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__9998 (
            .O(N__44617),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__9997 (
            .O(N__44610),
            .I(N__44607));
    LocalMux I__9996 (
            .O(N__44607),
            .I(N__44604));
    Span4Mux_v I__9995 (
            .O(N__44604),
            .I(N__44601));
    Odrv4 I__9994 (
            .O(N__44601),
            .I(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ));
    CascadeMux I__9993 (
            .O(N__44598),
            .I(N__44577));
    CascadeMux I__9992 (
            .O(N__44597),
            .I(N__44571));
    CascadeMux I__9991 (
            .O(N__44596),
            .I(N__44566));
    InMux I__9990 (
            .O(N__44595),
            .I(N__44560));
    InMux I__9989 (
            .O(N__44594),
            .I(N__44560));
    CascadeMux I__9988 (
            .O(N__44593),
            .I(N__44556));
    CascadeMux I__9987 (
            .O(N__44592),
            .I(N__44551));
    CascadeMux I__9986 (
            .O(N__44591),
            .I(N__44548));
    CascadeMux I__9985 (
            .O(N__44590),
            .I(N__44545));
    InMux I__9984 (
            .O(N__44589),
            .I(N__44542));
    InMux I__9983 (
            .O(N__44588),
            .I(N__44539));
    InMux I__9982 (
            .O(N__44587),
            .I(N__44536));
    InMux I__9981 (
            .O(N__44586),
            .I(N__44532));
    CascadeMux I__9980 (
            .O(N__44585),
            .I(N__44528));
    CascadeMux I__9979 (
            .O(N__44584),
            .I(N__44525));
    CascadeMux I__9978 (
            .O(N__44583),
            .I(N__44519));
    InMux I__9977 (
            .O(N__44582),
            .I(N__44505));
    InMux I__9976 (
            .O(N__44581),
            .I(N__44505));
    InMux I__9975 (
            .O(N__44580),
            .I(N__44502));
    InMux I__9974 (
            .O(N__44577),
            .I(N__44499));
    InMux I__9973 (
            .O(N__44576),
            .I(N__44496));
    InMux I__9972 (
            .O(N__44575),
            .I(N__44492));
    InMux I__9971 (
            .O(N__44574),
            .I(N__44481));
    InMux I__9970 (
            .O(N__44571),
            .I(N__44481));
    InMux I__9969 (
            .O(N__44570),
            .I(N__44481));
    InMux I__9968 (
            .O(N__44569),
            .I(N__44481));
    InMux I__9967 (
            .O(N__44566),
            .I(N__44481));
    InMux I__9966 (
            .O(N__44565),
            .I(N__44478));
    LocalMux I__9965 (
            .O(N__44560),
            .I(N__44475));
    InMux I__9964 (
            .O(N__44559),
            .I(N__44461));
    InMux I__9963 (
            .O(N__44556),
            .I(N__44461));
    InMux I__9962 (
            .O(N__44555),
            .I(N__44461));
    InMux I__9961 (
            .O(N__44554),
            .I(N__44461));
    InMux I__9960 (
            .O(N__44551),
            .I(N__44461));
    InMux I__9959 (
            .O(N__44548),
            .I(N__44461));
    InMux I__9958 (
            .O(N__44545),
            .I(N__44458));
    LocalMux I__9957 (
            .O(N__44542),
            .I(N__44453));
    LocalMux I__9956 (
            .O(N__44539),
            .I(N__44453));
    LocalMux I__9955 (
            .O(N__44536),
            .I(N__44450));
    InMux I__9954 (
            .O(N__44535),
            .I(N__44447));
    LocalMux I__9953 (
            .O(N__44532),
            .I(N__44444));
    InMux I__9952 (
            .O(N__44531),
            .I(N__44427));
    InMux I__9951 (
            .O(N__44528),
            .I(N__44427));
    InMux I__9950 (
            .O(N__44525),
            .I(N__44427));
    InMux I__9949 (
            .O(N__44524),
            .I(N__44427));
    InMux I__9948 (
            .O(N__44523),
            .I(N__44427));
    InMux I__9947 (
            .O(N__44522),
            .I(N__44427));
    InMux I__9946 (
            .O(N__44519),
            .I(N__44427));
    InMux I__9945 (
            .O(N__44518),
            .I(N__44427));
    InMux I__9944 (
            .O(N__44517),
            .I(N__44420));
    InMux I__9943 (
            .O(N__44516),
            .I(N__44420));
    InMux I__9942 (
            .O(N__44515),
            .I(N__44420));
    InMux I__9941 (
            .O(N__44514),
            .I(N__44417));
    InMux I__9940 (
            .O(N__44513),
            .I(N__44414));
    InMux I__9939 (
            .O(N__44512),
            .I(N__44407));
    InMux I__9938 (
            .O(N__44511),
            .I(N__44407));
    InMux I__9937 (
            .O(N__44510),
            .I(N__44407));
    LocalMux I__9936 (
            .O(N__44505),
            .I(N__44404));
    LocalMux I__9935 (
            .O(N__44502),
            .I(N__44401));
    LocalMux I__9934 (
            .O(N__44499),
            .I(N__44397));
    LocalMux I__9933 (
            .O(N__44496),
            .I(N__44394));
    InMux I__9932 (
            .O(N__44495),
            .I(N__44391));
    LocalMux I__9931 (
            .O(N__44492),
            .I(N__44386));
    LocalMux I__9930 (
            .O(N__44481),
            .I(N__44386));
    LocalMux I__9929 (
            .O(N__44478),
            .I(N__44381));
    Span4Mux_h I__9928 (
            .O(N__44475),
            .I(N__44381));
    CascadeMux I__9927 (
            .O(N__44474),
            .I(N__44377));
    LocalMux I__9926 (
            .O(N__44461),
            .I(N__44371));
    LocalMux I__9925 (
            .O(N__44458),
            .I(N__44368));
    Span4Mux_v I__9924 (
            .O(N__44453),
            .I(N__44365));
    Span4Mux_v I__9923 (
            .O(N__44450),
            .I(N__44358));
    LocalMux I__9922 (
            .O(N__44447),
            .I(N__44358));
    Span4Mux_h I__9921 (
            .O(N__44444),
            .I(N__44358));
    LocalMux I__9920 (
            .O(N__44427),
            .I(N__44353));
    LocalMux I__9919 (
            .O(N__44420),
            .I(N__44353));
    LocalMux I__9918 (
            .O(N__44417),
            .I(N__44342));
    LocalMux I__9917 (
            .O(N__44414),
            .I(N__44342));
    LocalMux I__9916 (
            .O(N__44407),
            .I(N__44342));
    Span4Mux_h I__9915 (
            .O(N__44404),
            .I(N__44342));
    Span4Mux_h I__9914 (
            .O(N__44401),
            .I(N__44342));
    InMux I__9913 (
            .O(N__44400),
            .I(N__44339));
    Span4Mux_h I__9912 (
            .O(N__44397),
            .I(N__44336));
    Span4Mux_h I__9911 (
            .O(N__44394),
            .I(N__44333));
    LocalMux I__9910 (
            .O(N__44391),
            .I(N__44330));
    Span4Mux_h I__9909 (
            .O(N__44386),
            .I(N__44325));
    Span4Mux_h I__9908 (
            .O(N__44381),
            .I(N__44325));
    InMux I__9907 (
            .O(N__44380),
            .I(N__44314));
    InMux I__9906 (
            .O(N__44377),
            .I(N__44314));
    InMux I__9905 (
            .O(N__44376),
            .I(N__44314));
    InMux I__9904 (
            .O(N__44375),
            .I(N__44314));
    InMux I__9903 (
            .O(N__44374),
            .I(N__44314));
    Span4Mux_h I__9902 (
            .O(N__44371),
            .I(N__44305));
    Span4Mux_h I__9901 (
            .O(N__44368),
            .I(N__44305));
    Span4Mux_h I__9900 (
            .O(N__44365),
            .I(N__44305));
    Span4Mux_v I__9899 (
            .O(N__44358),
            .I(N__44305));
    Span4Mux_h I__9898 (
            .O(N__44353),
            .I(N__44300));
    Span4Mux_v I__9897 (
            .O(N__44342),
            .I(N__44300));
    LocalMux I__9896 (
            .O(N__44339),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__9895 (
            .O(N__44336),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__9894 (
            .O(N__44333),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv12 I__9893 (
            .O(N__44330),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__9892 (
            .O(N__44325),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    LocalMux I__9891 (
            .O(N__44314),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__9890 (
            .O(N__44305),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__9889 (
            .O(N__44300),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__9888 (
            .O(N__44283),
            .I(N__44279));
    InMux I__9887 (
            .O(N__44282),
            .I(N__44276));
    LocalMux I__9886 (
            .O(N__44279),
            .I(N__44273));
    LocalMux I__9885 (
            .O(N__44276),
            .I(N__44270));
    Span4Mux_h I__9884 (
            .O(N__44273),
            .I(N__44266));
    Span4Mux_h I__9883 (
            .O(N__44270),
            .I(N__44263));
    InMux I__9882 (
            .O(N__44269),
            .I(N__44260));
    Span4Mux_h I__9881 (
            .O(N__44266),
            .I(N__44257));
    Span4Mux_h I__9880 (
            .O(N__44263),
            .I(N__44254));
    LocalMux I__9879 (
            .O(N__44260),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    Odrv4 I__9878 (
            .O(N__44257),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    Odrv4 I__9877 (
            .O(N__44254),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    InMux I__9876 (
            .O(N__44247),
            .I(N__44244));
    LocalMux I__9875 (
            .O(N__44244),
            .I(N__44240));
    CascadeMux I__9874 (
            .O(N__44243),
            .I(N__44237));
    Span4Mux_v I__9873 (
            .O(N__44240),
            .I(N__44233));
    InMux I__9872 (
            .O(N__44237),
            .I(N__44230));
    InMux I__9871 (
            .O(N__44236),
            .I(N__44227));
    Odrv4 I__9870 (
            .O(N__44233),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__9869 (
            .O(N__44230),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__9868 (
            .O(N__44227),
            .I(\current_shift_inst.un4_control_input1_19 ));
    CascadeMux I__9867 (
            .O(N__44220),
            .I(N__44217));
    InMux I__9866 (
            .O(N__44217),
            .I(N__44213));
    InMux I__9865 (
            .O(N__44216),
            .I(N__44209));
    LocalMux I__9864 (
            .O(N__44213),
            .I(N__44206));
    InMux I__9863 (
            .O(N__44212),
            .I(N__44203));
    LocalMux I__9862 (
            .O(N__44209),
            .I(N__44200));
    Span4Mux_v I__9861 (
            .O(N__44206),
            .I(N__44194));
    LocalMux I__9860 (
            .O(N__44203),
            .I(N__44194));
    Span4Mux_v I__9859 (
            .O(N__44200),
            .I(N__44191));
    InMux I__9858 (
            .O(N__44199),
            .I(N__44188));
    Sp12to4 I__9857 (
            .O(N__44194),
            .I(N__44181));
    Sp12to4 I__9856 (
            .O(N__44191),
            .I(N__44181));
    LocalMux I__9855 (
            .O(N__44188),
            .I(N__44181));
    Odrv12 I__9854 (
            .O(N__44181),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    CascadeMux I__9853 (
            .O(N__44178),
            .I(N__44175));
    InMux I__9852 (
            .O(N__44175),
            .I(N__44172));
    LocalMux I__9851 (
            .O(N__44172),
            .I(N__44169));
    Span4Mux_v I__9850 (
            .O(N__44169),
            .I(N__44166));
    Odrv4 I__9849 (
            .O(N__44166),
            .I(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ));
    InMux I__9848 (
            .O(N__44163),
            .I(N__44160));
    LocalMux I__9847 (
            .O(N__44160),
            .I(N__44156));
    InMux I__9846 (
            .O(N__44159),
            .I(N__44152));
    Span4Mux_v I__9845 (
            .O(N__44156),
            .I(N__44149));
    InMux I__9844 (
            .O(N__44155),
            .I(N__44146));
    LocalMux I__9843 (
            .O(N__44152),
            .I(N__44143));
    Odrv4 I__9842 (
            .O(N__44149),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__9841 (
            .O(N__44146),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__9840 (
            .O(N__44143),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    CEMux I__9839 (
            .O(N__44136),
            .I(N__44109));
    CEMux I__9838 (
            .O(N__44135),
            .I(N__44109));
    CEMux I__9837 (
            .O(N__44134),
            .I(N__44109));
    CEMux I__9836 (
            .O(N__44133),
            .I(N__44109));
    CEMux I__9835 (
            .O(N__44132),
            .I(N__44109));
    CEMux I__9834 (
            .O(N__44131),
            .I(N__44109));
    CEMux I__9833 (
            .O(N__44130),
            .I(N__44109));
    CEMux I__9832 (
            .O(N__44129),
            .I(N__44109));
    CEMux I__9831 (
            .O(N__44128),
            .I(N__44109));
    GlobalMux I__9830 (
            .O(N__44109),
            .I(N__44106));
    gio2CtrlBuf I__9829 (
            .O(N__44106),
            .I(\current_shift_inst.timer_s1.N_166_i_g ));
    CascadeMux I__9828 (
            .O(N__44103),
            .I(N__44099));
    InMux I__9827 (
            .O(N__44102),
            .I(N__44094));
    InMux I__9826 (
            .O(N__44099),
            .I(N__44094));
    LocalMux I__9825 (
            .O(N__44094),
            .I(N__44090));
    InMux I__9824 (
            .O(N__44093),
            .I(N__44087));
    Span4Mux_h I__9823 (
            .O(N__44090),
            .I(N__44081));
    LocalMux I__9822 (
            .O(N__44087),
            .I(N__44081));
    InMux I__9821 (
            .O(N__44086),
            .I(N__44078));
    Span4Mux_v I__9820 (
            .O(N__44081),
            .I(N__44075));
    LocalMux I__9819 (
            .O(N__44078),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__9818 (
            .O(N__44075),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__9817 (
            .O(N__44070),
            .I(N__44067));
    InMux I__9816 (
            .O(N__44067),
            .I(N__44064));
    LocalMux I__9815 (
            .O(N__44064),
            .I(N__44061));
    Span4Mux_h I__9814 (
            .O(N__44061),
            .I(N__44058));
    Odrv4 I__9813 (
            .O(N__44058),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__9812 (
            .O(N__44055),
            .I(N__44042));
    InMux I__9811 (
            .O(N__44054),
            .I(N__44033));
    InMux I__9810 (
            .O(N__44053),
            .I(N__44028));
    InMux I__9809 (
            .O(N__44052),
            .I(N__44028));
    InMux I__9808 (
            .O(N__44051),
            .I(N__44025));
    InMux I__9807 (
            .O(N__44050),
            .I(N__44004));
    InMux I__9806 (
            .O(N__44049),
            .I(N__44004));
    InMux I__9805 (
            .O(N__44048),
            .I(N__44004));
    InMux I__9804 (
            .O(N__44047),
            .I(N__44004));
    InMux I__9803 (
            .O(N__44046),
            .I(N__44004));
    InMux I__9802 (
            .O(N__44045),
            .I(N__44004));
    LocalMux I__9801 (
            .O(N__44042),
            .I(N__44001));
    InMux I__9800 (
            .O(N__44041),
            .I(N__43992));
    InMux I__9799 (
            .O(N__44040),
            .I(N__43992));
    InMux I__9798 (
            .O(N__44039),
            .I(N__43992));
    InMux I__9797 (
            .O(N__44038),
            .I(N__43992));
    InMux I__9796 (
            .O(N__44037),
            .I(N__43987));
    InMux I__9795 (
            .O(N__44036),
            .I(N__43987));
    LocalMux I__9794 (
            .O(N__44033),
            .I(N__43984));
    LocalMux I__9793 (
            .O(N__44028),
            .I(N__43981));
    LocalMux I__9792 (
            .O(N__44025),
            .I(N__43978));
    InMux I__9791 (
            .O(N__44024),
            .I(N__43975));
    InMux I__9790 (
            .O(N__44023),
            .I(N__43960));
    InMux I__9789 (
            .O(N__44022),
            .I(N__43960));
    InMux I__9788 (
            .O(N__44021),
            .I(N__43960));
    InMux I__9787 (
            .O(N__44020),
            .I(N__43960));
    InMux I__9786 (
            .O(N__44019),
            .I(N__43960));
    InMux I__9785 (
            .O(N__44018),
            .I(N__43960));
    InMux I__9784 (
            .O(N__44017),
            .I(N__43960));
    LocalMux I__9783 (
            .O(N__44004),
            .I(N__43955));
    Span4Mux_h I__9782 (
            .O(N__44001),
            .I(N__43955));
    LocalMux I__9781 (
            .O(N__43992),
            .I(N__43952));
    LocalMux I__9780 (
            .O(N__43987),
            .I(N__43945));
    Span4Mux_v I__9779 (
            .O(N__43984),
            .I(N__43945));
    Span4Mux_v I__9778 (
            .O(N__43981),
            .I(N__43945));
    Odrv4 I__9777 (
            .O(N__43978),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__9776 (
            .O(N__43975),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__9775 (
            .O(N__43960),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__9774 (
            .O(N__43955),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv12 I__9773 (
            .O(N__43952),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__9772 (
            .O(N__43945),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    CascadeMux I__9771 (
            .O(N__43932),
            .I(N__43928));
    InMux I__9770 (
            .O(N__43931),
            .I(N__43920));
    InMux I__9769 (
            .O(N__43928),
            .I(N__43920));
    InMux I__9768 (
            .O(N__43927),
            .I(N__43920));
    LocalMux I__9767 (
            .O(N__43920),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__9766 (
            .O(N__43917),
            .I(N__43907));
    InMux I__9765 (
            .O(N__43916),
            .I(N__43907));
    InMux I__9764 (
            .O(N__43915),
            .I(N__43907));
    InMux I__9763 (
            .O(N__43914),
            .I(N__43904));
    LocalMux I__9762 (
            .O(N__43907),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__9761 (
            .O(N__43904),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__9760 (
            .O(N__43899),
            .I(N__43896));
    InMux I__9759 (
            .O(N__43896),
            .I(N__43893));
    LocalMux I__9758 (
            .O(N__43893),
            .I(N__43890));
    Span4Mux_h I__9757 (
            .O(N__43890),
            .I(N__43887));
    Odrv4 I__9756 (
            .O(N__43887),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    CascadeMux I__9755 (
            .O(N__43884),
            .I(N__43881));
    InMux I__9754 (
            .O(N__43881),
            .I(N__43878));
    LocalMux I__9753 (
            .O(N__43878),
            .I(N__43875));
    Span4Mux_h I__9752 (
            .O(N__43875),
            .I(N__43872));
    Odrv4 I__9751 (
            .O(N__43872),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    CascadeMux I__9750 (
            .O(N__43869),
            .I(N__43866));
    InMux I__9749 (
            .O(N__43866),
            .I(N__43863));
    LocalMux I__9748 (
            .O(N__43863),
            .I(N__43860));
    Span12Mux_h I__9747 (
            .O(N__43860),
            .I(N__43857));
    Odrv12 I__9746 (
            .O(N__43857),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    CascadeMux I__9745 (
            .O(N__43854),
            .I(N__43851));
    InMux I__9744 (
            .O(N__43851),
            .I(N__43847));
    InMux I__9743 (
            .O(N__43850),
            .I(N__43844));
    LocalMux I__9742 (
            .O(N__43847),
            .I(N__43836));
    LocalMux I__9741 (
            .O(N__43844),
            .I(N__43836));
    InMux I__9740 (
            .O(N__43843),
            .I(N__43831));
    InMux I__9739 (
            .O(N__43842),
            .I(N__43831));
    InMux I__9738 (
            .O(N__43841),
            .I(N__43828));
    Span4Mux_h I__9737 (
            .O(N__43836),
            .I(N__43823));
    LocalMux I__9736 (
            .O(N__43831),
            .I(N__43823));
    LocalMux I__9735 (
            .O(N__43828),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__9734 (
            .O(N__43823),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__9733 (
            .O(N__43818),
            .I(N__43813));
    InMux I__9732 (
            .O(N__43817),
            .I(N__43808));
    InMux I__9731 (
            .O(N__43816),
            .I(N__43808));
    LocalMux I__9730 (
            .O(N__43813),
            .I(N__43803));
    LocalMux I__9729 (
            .O(N__43808),
            .I(N__43803));
    Odrv4 I__9728 (
            .O(N__43803),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__9727 (
            .O(N__43800),
            .I(N__43797));
    InMux I__9726 (
            .O(N__43797),
            .I(N__43794));
    LocalMux I__9725 (
            .O(N__43794),
            .I(N__43791));
    Span4Mux_h I__9724 (
            .O(N__43791),
            .I(N__43788));
    Span4Mux_v I__9723 (
            .O(N__43788),
            .I(N__43785));
    Odrv4 I__9722 (
            .O(N__43785),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    CascadeMux I__9721 (
            .O(N__43782),
            .I(N__43779));
    InMux I__9720 (
            .O(N__43779),
            .I(N__43776));
    LocalMux I__9719 (
            .O(N__43776),
            .I(N__43770));
    InMux I__9718 (
            .O(N__43775),
            .I(N__43765));
    InMux I__9717 (
            .O(N__43774),
            .I(N__43765));
    InMux I__9716 (
            .O(N__43773),
            .I(N__43762));
    Span4Mux_v I__9715 (
            .O(N__43770),
            .I(N__43759));
    LocalMux I__9714 (
            .O(N__43765),
            .I(N__43756));
    LocalMux I__9713 (
            .O(N__43762),
            .I(N__43753));
    Span4Mux_h I__9712 (
            .O(N__43759),
            .I(N__43750));
    Span4Mux_h I__9711 (
            .O(N__43756),
            .I(N__43747));
    Odrv4 I__9710 (
            .O(N__43753),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__9709 (
            .O(N__43750),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__9708 (
            .O(N__43747),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    CascadeMux I__9707 (
            .O(N__43740),
            .I(N__43737));
    InMux I__9706 (
            .O(N__43737),
            .I(N__43733));
    InMux I__9705 (
            .O(N__43736),
            .I(N__43729));
    LocalMux I__9704 (
            .O(N__43733),
            .I(N__43726));
    InMux I__9703 (
            .O(N__43732),
            .I(N__43723));
    LocalMux I__9702 (
            .O(N__43729),
            .I(N__43718));
    Span4Mux_v I__9701 (
            .O(N__43726),
            .I(N__43718));
    LocalMux I__9700 (
            .O(N__43723),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__9699 (
            .O(N__43718),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__9698 (
            .O(N__43713),
            .I(N__43710));
    LocalMux I__9697 (
            .O(N__43710),
            .I(N__43707));
    Span4Mux_v I__9696 (
            .O(N__43707),
            .I(N__43704));
    Odrv4 I__9695 (
            .O(N__43704),
            .I(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ));
    CascadeMux I__9694 (
            .O(N__43701),
            .I(N__43697));
    CascadeMux I__9693 (
            .O(N__43700),
            .I(N__43694));
    InMux I__9692 (
            .O(N__43697),
            .I(N__43690));
    InMux I__9691 (
            .O(N__43694),
            .I(N__43687));
    InMux I__9690 (
            .O(N__43693),
            .I(N__43684));
    LocalMux I__9689 (
            .O(N__43690),
            .I(N__43680));
    LocalMux I__9688 (
            .O(N__43687),
            .I(N__43677));
    LocalMux I__9687 (
            .O(N__43684),
            .I(N__43674));
    InMux I__9686 (
            .O(N__43683),
            .I(N__43671));
    Span4Mux_h I__9685 (
            .O(N__43680),
            .I(N__43668));
    Span4Mux_v I__9684 (
            .O(N__43677),
            .I(N__43663));
    Span4Mux_h I__9683 (
            .O(N__43674),
            .I(N__43663));
    LocalMux I__9682 (
            .O(N__43671),
            .I(N__43660));
    Span4Mux_h I__9681 (
            .O(N__43668),
            .I(N__43657));
    Span4Mux_h I__9680 (
            .O(N__43663),
            .I(N__43654));
    Odrv12 I__9679 (
            .O(N__43660),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__9678 (
            .O(N__43657),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__9677 (
            .O(N__43654),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__9676 (
            .O(N__43647),
            .I(N__43643));
    InMux I__9675 (
            .O(N__43646),
            .I(N__43639));
    LocalMux I__9674 (
            .O(N__43643),
            .I(N__43636));
    InMux I__9673 (
            .O(N__43642),
            .I(N__43633));
    LocalMux I__9672 (
            .O(N__43639),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__9671 (
            .O(N__43636),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__9670 (
            .O(N__43633),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__9669 (
            .O(N__43626),
            .I(N__43623));
    InMux I__9668 (
            .O(N__43623),
            .I(N__43620));
    LocalMux I__9667 (
            .O(N__43620),
            .I(N__43617));
    Span4Mux_v I__9666 (
            .O(N__43617),
            .I(N__43614));
    Odrv4 I__9665 (
            .O(N__43614),
            .I(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ));
    InMux I__9664 (
            .O(N__43611),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__9663 (
            .O(N__43608),
            .I(N__43604));
    InMux I__9662 (
            .O(N__43607),
            .I(N__43600));
    InMux I__9661 (
            .O(N__43604),
            .I(N__43597));
    InMux I__9660 (
            .O(N__43603),
            .I(N__43594));
    LocalMux I__9659 (
            .O(N__43600),
            .I(N__43591));
    LocalMux I__9658 (
            .O(N__43597),
            .I(N__43588));
    LocalMux I__9657 (
            .O(N__43594),
            .I(N__43585));
    Span4Mux_v I__9656 (
            .O(N__43591),
            .I(N__43580));
    Span4Mux_h I__9655 (
            .O(N__43588),
            .I(N__43580));
    Span12Mux_h I__9654 (
            .O(N__43585),
            .I(N__43576));
    Span4Mux_h I__9653 (
            .O(N__43580),
            .I(N__43573));
    InMux I__9652 (
            .O(N__43579),
            .I(N__43570));
    Odrv12 I__9651 (
            .O(N__43576),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__9650 (
            .O(N__43573),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__9649 (
            .O(N__43570),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    CascadeMux I__9648 (
            .O(N__43563),
            .I(N__43560));
    InMux I__9647 (
            .O(N__43560),
            .I(N__43557));
    LocalMux I__9646 (
            .O(N__43557),
            .I(N__43554));
    Span4Mux_v I__9645 (
            .O(N__43554),
            .I(N__43549));
    InMux I__9644 (
            .O(N__43553),
            .I(N__43546));
    InMux I__9643 (
            .O(N__43552),
            .I(N__43543));
    Odrv4 I__9642 (
            .O(N__43549),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__9641 (
            .O(N__43546),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__9640 (
            .O(N__43543),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__9639 (
            .O(N__43536),
            .I(N__43533));
    InMux I__9638 (
            .O(N__43533),
            .I(N__43530));
    LocalMux I__9637 (
            .O(N__43530),
            .I(N__43527));
    Sp12to4 I__9636 (
            .O(N__43527),
            .I(N__43524));
    Odrv12 I__9635 (
            .O(N__43524),
            .I(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ));
    CascadeMux I__9634 (
            .O(N__43521),
            .I(N__43518));
    InMux I__9633 (
            .O(N__43518),
            .I(N__43515));
    LocalMux I__9632 (
            .O(N__43515),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__9631 (
            .O(N__43512),
            .I(N__43509));
    LocalMux I__9630 (
            .O(N__43509),
            .I(N__43506));
    Odrv4 I__9629 (
            .O(N__43506),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__9628 (
            .O(N__43503),
            .I(N__43499));
    CascadeMux I__9627 (
            .O(N__43502),
            .I(N__43496));
    InMux I__9626 (
            .O(N__43499),
            .I(N__43493));
    InMux I__9625 (
            .O(N__43496),
            .I(N__43490));
    LocalMux I__9624 (
            .O(N__43493),
            .I(N__43485));
    LocalMux I__9623 (
            .O(N__43490),
            .I(N__43482));
    InMux I__9622 (
            .O(N__43489),
            .I(N__43477));
    InMux I__9621 (
            .O(N__43488),
            .I(N__43477));
    Span4Mux_v I__9620 (
            .O(N__43485),
            .I(N__43474));
    Span12Mux_s7_v I__9619 (
            .O(N__43482),
            .I(N__43469));
    LocalMux I__9618 (
            .O(N__43477),
            .I(N__43469));
    Odrv4 I__9617 (
            .O(N__43474),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv12 I__9616 (
            .O(N__43469),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__9615 (
            .O(N__43464),
            .I(N__43461));
    LocalMux I__9614 (
            .O(N__43461),
            .I(N__43458));
    Span4Mux_v I__9613 (
            .O(N__43458),
            .I(N__43453));
    InMux I__9612 (
            .O(N__43457),
            .I(N__43450));
    InMux I__9611 (
            .O(N__43456),
            .I(N__43447));
    Odrv4 I__9610 (
            .O(N__43453),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__9609 (
            .O(N__43450),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__9608 (
            .O(N__43447),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__9607 (
            .O(N__43440),
            .I(N__43437));
    LocalMux I__9606 (
            .O(N__43437),
            .I(N__43434));
    Span4Mux_v I__9605 (
            .O(N__43434),
            .I(N__43431));
    Odrv4 I__9604 (
            .O(N__43431),
            .I(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ));
    CascadeMux I__9603 (
            .O(N__43428),
            .I(N__43425));
    InMux I__9602 (
            .O(N__43425),
            .I(N__43422));
    LocalMux I__9601 (
            .O(N__43422),
            .I(N__43418));
    CascadeMux I__9600 (
            .O(N__43421),
            .I(N__43415));
    Span4Mux_v I__9599 (
            .O(N__43418),
            .I(N__43410));
    InMux I__9598 (
            .O(N__43415),
            .I(N__43407));
    InMux I__9597 (
            .O(N__43414),
            .I(N__43402));
    InMux I__9596 (
            .O(N__43413),
            .I(N__43402));
    Span4Mux_h I__9595 (
            .O(N__43410),
            .I(N__43399));
    LocalMux I__9594 (
            .O(N__43407),
            .I(N__43396));
    LocalMux I__9593 (
            .O(N__43402),
            .I(N__43393));
    Odrv4 I__9592 (
            .O(N__43399),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv12 I__9591 (
            .O(N__43396),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__9590 (
            .O(N__43393),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__9589 (
            .O(N__43386),
            .I(N__43382));
    InMux I__9588 (
            .O(N__43385),
            .I(N__43379));
    LocalMux I__9587 (
            .O(N__43382),
            .I(N__43375));
    LocalMux I__9586 (
            .O(N__43379),
            .I(N__43372));
    InMux I__9585 (
            .O(N__43378),
            .I(N__43369));
    Span4Mux_v I__9584 (
            .O(N__43375),
            .I(N__43364));
    Span4Mux_h I__9583 (
            .O(N__43372),
            .I(N__43364));
    LocalMux I__9582 (
            .O(N__43369),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__9581 (
            .O(N__43364),
            .I(\current_shift_inst.un4_control_input1_7 ));
    CascadeMux I__9580 (
            .O(N__43359),
            .I(N__43356));
    InMux I__9579 (
            .O(N__43356),
            .I(N__43353));
    LocalMux I__9578 (
            .O(N__43353),
            .I(N__43350));
    Span4Mux_v I__9577 (
            .O(N__43350),
            .I(N__43347));
    Odrv4 I__9576 (
            .O(N__43347),
            .I(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ));
    InMux I__9575 (
            .O(N__43344),
            .I(N__43341));
    LocalMux I__9574 (
            .O(N__43341),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    CascadeMux I__9573 (
            .O(N__43338),
            .I(N__43335));
    InMux I__9572 (
            .O(N__43335),
            .I(N__43331));
    InMux I__9571 (
            .O(N__43334),
            .I(N__43328));
    LocalMux I__9570 (
            .O(N__43331),
            .I(N__43322));
    LocalMux I__9569 (
            .O(N__43328),
            .I(N__43322));
    InMux I__9568 (
            .O(N__43327),
            .I(N__43319));
    Odrv4 I__9567 (
            .O(N__43322),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__9566 (
            .O(N__43319),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__9565 (
            .O(N__43314),
            .I(N__43309));
    InMux I__9564 (
            .O(N__43313),
            .I(N__43306));
    CascadeMux I__9563 (
            .O(N__43312),
            .I(N__43303));
    LocalMux I__9562 (
            .O(N__43309),
            .I(N__43299));
    LocalMux I__9561 (
            .O(N__43306),
            .I(N__43296));
    InMux I__9560 (
            .O(N__43303),
            .I(N__43291));
    InMux I__9559 (
            .O(N__43302),
            .I(N__43291));
    Span4Mux_h I__9558 (
            .O(N__43299),
            .I(N__43284));
    Span4Mux_v I__9557 (
            .O(N__43296),
            .I(N__43284));
    LocalMux I__9556 (
            .O(N__43291),
            .I(N__43284));
    Odrv4 I__9555 (
            .O(N__43284),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    CascadeMux I__9554 (
            .O(N__43281),
            .I(N__43278));
    InMux I__9553 (
            .O(N__43278),
            .I(N__43275));
    LocalMux I__9552 (
            .O(N__43275),
            .I(N__43272));
    Sp12to4 I__9551 (
            .O(N__43272),
            .I(N__43269));
    Odrv12 I__9550 (
            .O(N__43269),
            .I(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ));
    CascadeMux I__9549 (
            .O(N__43266),
            .I(N__43263));
    InMux I__9548 (
            .O(N__43263),
            .I(N__43260));
    LocalMux I__9547 (
            .O(N__43260),
            .I(N__43257));
    Span4Mux_h I__9546 (
            .O(N__43257),
            .I(N__43254));
    Span4Mux_v I__9545 (
            .O(N__43254),
            .I(N__43251));
    Odrv4 I__9544 (
            .O(N__43251),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ));
    CascadeMux I__9543 (
            .O(N__43248),
            .I(N__43245));
    InMux I__9542 (
            .O(N__43245),
            .I(N__43242));
    LocalMux I__9541 (
            .O(N__43242),
            .I(N__43238));
    InMux I__9540 (
            .O(N__43241),
            .I(N__43235));
    Odrv12 I__9539 (
            .O(N__43238),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__9538 (
            .O(N__43235),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__9537 (
            .O(N__43230),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__9536 (
            .O(N__43227),
            .I(N__43224));
    InMux I__9535 (
            .O(N__43224),
            .I(N__43221));
    LocalMux I__9534 (
            .O(N__43221),
            .I(N__43217));
    InMux I__9533 (
            .O(N__43220),
            .I(N__43214));
    Span4Mux_v I__9532 (
            .O(N__43217),
            .I(N__43209));
    LocalMux I__9531 (
            .O(N__43214),
            .I(N__43209));
    Odrv4 I__9530 (
            .O(N__43209),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__9529 (
            .O(N__43206),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__9528 (
            .O(N__43203),
            .I(N__43200));
    InMux I__9527 (
            .O(N__43200),
            .I(N__43196));
    CascadeMux I__9526 (
            .O(N__43199),
            .I(N__43193));
    LocalMux I__9525 (
            .O(N__43196),
            .I(N__43190));
    InMux I__9524 (
            .O(N__43193),
            .I(N__43187));
    Span4Mux_v I__9523 (
            .O(N__43190),
            .I(N__43182));
    LocalMux I__9522 (
            .O(N__43187),
            .I(N__43182));
    Odrv4 I__9521 (
            .O(N__43182),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__9520 (
            .O(N__43179),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__9519 (
            .O(N__43176),
            .I(N__43173));
    LocalMux I__9518 (
            .O(N__43173),
            .I(N__43170));
    Span4Mux_v I__9517 (
            .O(N__43170),
            .I(N__43166));
    InMux I__9516 (
            .O(N__43169),
            .I(N__43163));
    Odrv4 I__9515 (
            .O(N__43166),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    LocalMux I__9514 (
            .O(N__43163),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__9513 (
            .O(N__43158),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__9512 (
            .O(N__43155),
            .I(N__43152));
    LocalMux I__9511 (
            .O(N__43152),
            .I(N__43148));
    CascadeMux I__9510 (
            .O(N__43151),
            .I(N__43145));
    Span4Mux_v I__9509 (
            .O(N__43148),
            .I(N__43142));
    InMux I__9508 (
            .O(N__43145),
            .I(N__43139));
    Odrv4 I__9507 (
            .O(N__43142),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    LocalMux I__9506 (
            .O(N__43139),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__9505 (
            .O(N__43134),
            .I(bfn_17_22_0_));
    InMux I__9504 (
            .O(N__43131),
            .I(N__43128));
    LocalMux I__9503 (
            .O(N__43128),
            .I(N__43125));
    Span4Mux_v I__9502 (
            .O(N__43125),
            .I(N__43121));
    InMux I__9501 (
            .O(N__43124),
            .I(N__43118));
    Odrv4 I__9500 (
            .O(N__43121),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    LocalMux I__9499 (
            .O(N__43118),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__9498 (
            .O(N__43113),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__9497 (
            .O(N__43110),
            .I(N__43106));
    InMux I__9496 (
            .O(N__43109),
            .I(N__43103));
    LocalMux I__9495 (
            .O(N__43106),
            .I(N__43100));
    LocalMux I__9494 (
            .O(N__43103),
            .I(N__43097));
    Odrv12 I__9493 (
            .O(N__43100),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__9492 (
            .O(N__43097),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__9491 (
            .O(N__43092),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__9490 (
            .O(N__43089),
            .I(N__43085));
    InMux I__9489 (
            .O(N__43088),
            .I(N__43082));
    LocalMux I__9488 (
            .O(N__43085),
            .I(N__43079));
    LocalMux I__9487 (
            .O(N__43082),
            .I(N__43076));
    Odrv12 I__9486 (
            .O(N__43079),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__9485 (
            .O(N__43076),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__9484 (
            .O(N__43071),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__9483 (
            .O(N__43068),
            .I(N__43063));
    InMux I__9482 (
            .O(N__43067),
            .I(N__43057));
    InMux I__9481 (
            .O(N__43066),
            .I(N__43057));
    LocalMux I__9480 (
            .O(N__43063),
            .I(N__43054));
    InMux I__9479 (
            .O(N__43062),
            .I(N__43051));
    LocalMux I__9478 (
            .O(N__43057),
            .I(N__43048));
    Odrv4 I__9477 (
            .O(N__43054),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    LocalMux I__9476 (
            .O(N__43051),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    Odrv4 I__9475 (
            .O(N__43048),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    InMux I__9474 (
            .O(N__43041),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__9473 (
            .O(N__43038),
            .I(N__43034));
    InMux I__9472 (
            .O(N__43037),
            .I(N__43031));
    LocalMux I__9471 (
            .O(N__43034),
            .I(N__43028));
    LocalMux I__9470 (
            .O(N__43031),
            .I(N__43025));
    Span4Mux_v I__9469 (
            .O(N__43028),
            .I(N__43019));
    Span4Mux_h I__9468 (
            .O(N__43025),
            .I(N__43019));
    InMux I__9467 (
            .O(N__43024),
            .I(N__43016));
    Odrv4 I__9466 (
            .O(N__43019),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    LocalMux I__9465 (
            .O(N__43016),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    InMux I__9464 (
            .O(N__43011),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__9463 (
            .O(N__43008),
            .I(N__43003));
    CascadeMux I__9462 (
            .O(N__43007),
            .I(N__43000));
    CascadeMux I__9461 (
            .O(N__43006),
            .I(N__42997));
    LocalMux I__9460 (
            .O(N__43003),
            .I(N__42994));
    InMux I__9459 (
            .O(N__43000),
            .I(N__42991));
    InMux I__9458 (
            .O(N__42997),
            .I(N__42988));
    Odrv4 I__9457 (
            .O(N__42994),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__9456 (
            .O(N__42991),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__9455 (
            .O(N__42988),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__9454 (
            .O(N__42981),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__9453 (
            .O(N__42978),
            .I(N__42975));
    LocalMux I__9452 (
            .O(N__42975),
            .I(N__42971));
    InMux I__9451 (
            .O(N__42974),
            .I(N__42968));
    Span4Mux_v I__9450 (
            .O(N__42971),
            .I(N__42964));
    LocalMux I__9449 (
            .O(N__42968),
            .I(N__42961));
    InMux I__9448 (
            .O(N__42967),
            .I(N__42958));
    Odrv4 I__9447 (
            .O(N__42964),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv4 I__9446 (
            .O(N__42961),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__9445 (
            .O(N__42958),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__9444 (
            .O(N__42951),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__9443 (
            .O(N__42948),
            .I(N__42945));
    LocalMux I__9442 (
            .O(N__42945),
            .I(N__42942));
    Span4Mux_v I__9441 (
            .O(N__42942),
            .I(N__42937));
    InMux I__9440 (
            .O(N__42941),
            .I(N__42934));
    InMux I__9439 (
            .O(N__42940),
            .I(N__42931));
    Odrv4 I__9438 (
            .O(N__42937),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__9437 (
            .O(N__42934),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__9436 (
            .O(N__42931),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__9435 (
            .O(N__42924),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__9434 (
            .O(N__42921),
            .I(bfn_17_21_0_));
    CascadeMux I__9433 (
            .O(N__42918),
            .I(N__42915));
    InMux I__9432 (
            .O(N__42915),
            .I(N__42912));
    LocalMux I__9431 (
            .O(N__42912),
            .I(N__42909));
    Span4Mux_v I__9430 (
            .O(N__42909),
            .I(N__42905));
    InMux I__9429 (
            .O(N__42908),
            .I(N__42902));
    Odrv4 I__9428 (
            .O(N__42905),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__9427 (
            .O(N__42902),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__9426 (
            .O(N__42897),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__9425 (
            .O(N__42894),
            .I(N__42891));
    LocalMux I__9424 (
            .O(N__42891),
            .I(N__42886));
    InMux I__9423 (
            .O(N__42890),
            .I(N__42881));
    InMux I__9422 (
            .O(N__42889),
            .I(N__42881));
    Span4Mux_v I__9421 (
            .O(N__42886),
            .I(N__42876));
    LocalMux I__9420 (
            .O(N__42881),
            .I(N__42876));
    Odrv4 I__9419 (
            .O(N__42876),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__9418 (
            .O(N__42873),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__9417 (
            .O(N__42870),
            .I(N__42865));
    InMux I__9416 (
            .O(N__42869),
            .I(N__42860));
    InMux I__9415 (
            .O(N__42868),
            .I(N__42860));
    LocalMux I__9414 (
            .O(N__42865),
            .I(N__42857));
    LocalMux I__9413 (
            .O(N__42860),
            .I(N__42854));
    Span4Mux_v I__9412 (
            .O(N__42857),
            .I(N__42849));
    Span4Mux_h I__9411 (
            .O(N__42854),
            .I(N__42849));
    Odrv4 I__9410 (
            .O(N__42849),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__9409 (
            .O(N__42846),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__9408 (
            .O(N__42843),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__9407 (
            .O(N__42840),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__9406 (
            .O(N__42837),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__9405 (
            .O(N__42834),
            .I(N__42831));
    LocalMux I__9404 (
            .O(N__42831),
            .I(N__42826));
    CascadeMux I__9403 (
            .O(N__42830),
            .I(N__42822));
    CascadeMux I__9402 (
            .O(N__42829),
            .I(N__42819));
    Span4Mux_h I__9401 (
            .O(N__42826),
            .I(N__42816));
    InMux I__9400 (
            .O(N__42825),
            .I(N__42813));
    InMux I__9399 (
            .O(N__42822),
            .I(N__42810));
    InMux I__9398 (
            .O(N__42819),
            .I(N__42807));
    Odrv4 I__9397 (
            .O(N__42816),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    LocalMux I__9396 (
            .O(N__42813),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    LocalMux I__9395 (
            .O(N__42810),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    LocalMux I__9394 (
            .O(N__42807),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    InMux I__9393 (
            .O(N__42798),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__9392 (
            .O(N__42795),
            .I(N__42792));
    LocalMux I__9391 (
            .O(N__42792),
            .I(N__42788));
    InMux I__9390 (
            .O(N__42791),
            .I(N__42785));
    Odrv12 I__9389 (
            .O(N__42788),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__9388 (
            .O(N__42785),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__9387 (
            .O(N__42780),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__9386 (
            .O(N__42777),
            .I(N__42774));
    LocalMux I__9385 (
            .O(N__42774),
            .I(N__42770));
    InMux I__9384 (
            .O(N__42773),
            .I(N__42767));
    Odrv12 I__9383 (
            .O(N__42770),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__9382 (
            .O(N__42767),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__9381 (
            .O(N__42762),
            .I(bfn_17_20_0_));
    InMux I__9380 (
            .O(N__42759),
            .I(N__42756));
    LocalMux I__9379 (
            .O(N__42756),
            .I(N__42752));
    CascadeMux I__9378 (
            .O(N__42755),
            .I(N__42749));
    Span4Mux_h I__9377 (
            .O(N__42752),
            .I(N__42746));
    InMux I__9376 (
            .O(N__42749),
            .I(N__42743));
    Odrv4 I__9375 (
            .O(N__42746),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    LocalMux I__9374 (
            .O(N__42743),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__9373 (
            .O(N__42738),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__9372 (
            .O(N__42735),
            .I(N__42732));
    LocalMux I__9371 (
            .O(N__42732),
            .I(N__42729));
    Span4Mux_v I__9370 (
            .O(N__42729),
            .I(N__42725));
    InMux I__9369 (
            .O(N__42728),
            .I(N__42722));
    Odrv4 I__9368 (
            .O(N__42725),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__9367 (
            .O(N__42722),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__9366 (
            .O(N__42717),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__9365 (
            .O(N__42714),
            .I(N__42711));
    LocalMux I__9364 (
            .O(N__42711),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4 ));
    CascadeMux I__9363 (
            .O(N__42708),
            .I(N__42705));
    InMux I__9362 (
            .O(N__42705),
            .I(N__42702));
    LocalMux I__9361 (
            .O(N__42702),
            .I(\delay_measurement_inst.delay_tr_timer.N_344 ));
    CascadeMux I__9360 (
            .O(N__42699),
            .I(\delay_measurement_inst.delay_tr_timer.N_344_cascade_ ));
    InMux I__9359 (
            .O(N__42696),
            .I(N__42693));
    LocalMux I__9358 (
            .O(N__42693),
            .I(\delay_measurement_inst.delay_tr_timer.N_347 ));
    CascadeMux I__9357 (
            .O(N__42690),
            .I(\delay_measurement_inst.delay_tr_timer.N_347_cascade_ ));
    CascadeMux I__9356 (
            .O(N__42687),
            .I(\delay_measurement_inst.delay_tr_timer.N_373_cascade_ ));
    InMux I__9355 (
            .O(N__42684),
            .I(N__42681));
    LocalMux I__9354 (
            .O(N__42681),
            .I(\delay_measurement_inst.delay_tr_timer.N_351 ));
    InMux I__9353 (
            .O(N__42678),
            .I(N__42675));
    LocalMux I__9352 (
            .O(N__42675),
            .I(\delay_measurement_inst.delay_tr_timer.N_353 ));
    InMux I__9351 (
            .O(N__42672),
            .I(N__42668));
    InMux I__9350 (
            .O(N__42671),
            .I(N__42665));
    LocalMux I__9349 (
            .O(N__42668),
            .I(\delay_measurement_inst.delay_tr_timer.N_348 ));
    LocalMux I__9348 (
            .O(N__42665),
            .I(\delay_measurement_inst.delay_tr_timer.N_348 ));
    CascadeMux I__9347 (
            .O(N__42660),
            .I(N__42657));
    InMux I__9346 (
            .O(N__42657),
            .I(N__42654));
    LocalMux I__9345 (
            .O(N__42654),
            .I(N__42649));
    InMux I__9344 (
            .O(N__42653),
            .I(N__42644));
    InMux I__9343 (
            .O(N__42652),
            .I(N__42644));
    Odrv12 I__9342 (
            .O(N__42649),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__9341 (
            .O(N__42644),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__9340 (
            .O(N__42639),
            .I(N__42636));
    LocalMux I__9339 (
            .O(N__42636),
            .I(N__42632));
    InMux I__9338 (
            .O(N__42635),
            .I(N__42629));
    Odrv4 I__9337 (
            .O(N__42632),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__9336 (
            .O(N__42629),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__9335 (
            .O(N__42624),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__9334 (
            .O(N__42621),
            .I(N__42618));
    LocalMux I__9333 (
            .O(N__42618),
            .I(N__42614));
    InMux I__9332 (
            .O(N__42617),
            .I(N__42611));
    Odrv4 I__9331 (
            .O(N__42614),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__9330 (
            .O(N__42611),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__9329 (
            .O(N__42606),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__9328 (
            .O(N__42603),
            .I(N__42600));
    InMux I__9327 (
            .O(N__42600),
            .I(N__42596));
    InMux I__9326 (
            .O(N__42599),
            .I(N__42593));
    LocalMux I__9325 (
            .O(N__42596),
            .I(elapsed_time_ns_1_RNI3JIF91_0_29));
    LocalMux I__9324 (
            .O(N__42593),
            .I(elapsed_time_ns_1_RNI3JIF91_0_29));
    InMux I__9323 (
            .O(N__42588),
            .I(N__42585));
    LocalMux I__9322 (
            .O(N__42585),
            .I(elapsed_time_ns_1_RNITCIF91_0_23));
    CascadeMux I__9321 (
            .O(N__42582),
            .I(elapsed_time_ns_1_RNITCIF91_0_23_cascade_));
    InMux I__9320 (
            .O(N__42579),
            .I(N__42575));
    InMux I__9319 (
            .O(N__42578),
            .I(N__42572));
    LocalMux I__9318 (
            .O(N__42575),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    LocalMux I__9317 (
            .O(N__42572),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    InMux I__9316 (
            .O(N__42567),
            .I(N__42564));
    LocalMux I__9315 (
            .O(N__42564),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ));
    InMux I__9314 (
            .O(N__42561),
            .I(N__42557));
    InMux I__9313 (
            .O(N__42560),
            .I(N__42551));
    LocalMux I__9312 (
            .O(N__42557),
            .I(N__42548));
    InMux I__9311 (
            .O(N__42556),
            .I(N__42545));
    InMux I__9310 (
            .O(N__42555),
            .I(N__42542));
    InMux I__9309 (
            .O(N__42554),
            .I(N__42539));
    LocalMux I__9308 (
            .O(N__42551),
            .I(elapsed_time_ns_1_RNIA965M1_0_18));
    Odrv12 I__9307 (
            .O(N__42548),
            .I(elapsed_time_ns_1_RNIA965M1_0_18));
    LocalMux I__9306 (
            .O(N__42545),
            .I(elapsed_time_ns_1_RNIA965M1_0_18));
    LocalMux I__9305 (
            .O(N__42542),
            .I(elapsed_time_ns_1_RNIA965M1_0_18));
    LocalMux I__9304 (
            .O(N__42539),
            .I(elapsed_time_ns_1_RNIA965M1_0_18));
    CascadeMux I__9303 (
            .O(N__42528),
            .I(elapsed_time_ns_1_RNICG2591_0_4_cascade_));
    InMux I__9302 (
            .O(N__42525),
            .I(N__42522));
    LocalMux I__9301 (
            .O(N__42522),
            .I(N__42518));
    InMux I__9300 (
            .O(N__42521),
            .I(N__42512));
    Span4Mux_v I__9299 (
            .O(N__42518),
            .I(N__42509));
    InMux I__9298 (
            .O(N__42517),
            .I(N__42506));
    InMux I__9297 (
            .O(N__42516),
            .I(N__42503));
    InMux I__9296 (
            .O(N__42515),
            .I(N__42500));
    LocalMux I__9295 (
            .O(N__42512),
            .I(elapsed_time_ns_1_RNI9865M1_0_17));
    Odrv4 I__9294 (
            .O(N__42509),
            .I(elapsed_time_ns_1_RNI9865M1_0_17));
    LocalMux I__9293 (
            .O(N__42506),
            .I(elapsed_time_ns_1_RNI9865M1_0_17));
    LocalMux I__9292 (
            .O(N__42503),
            .I(elapsed_time_ns_1_RNI9865M1_0_17));
    LocalMux I__9291 (
            .O(N__42500),
            .I(elapsed_time_ns_1_RNI9865M1_0_17));
    CascadeMux I__9290 (
            .O(N__42489),
            .I(N__42486));
    InMux I__9289 (
            .O(N__42486),
            .I(N__42482));
    InMux I__9288 (
            .O(N__42485),
            .I(N__42479));
    LocalMux I__9287 (
            .O(N__42482),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9 ));
    LocalMux I__9286 (
            .O(N__42479),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9 ));
    CascadeMux I__9285 (
            .O(N__42474),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_ ));
    CascadeMux I__9284 (
            .O(N__42471),
            .I(N__42468));
    InMux I__9283 (
            .O(N__42468),
            .I(N__42464));
    InMux I__9282 (
            .O(N__42467),
            .I(N__42461));
    LocalMux I__9281 (
            .O(N__42464),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    LocalMux I__9280 (
            .O(N__42461),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    InMux I__9279 (
            .O(N__42456),
            .I(N__42453));
    LocalMux I__9278 (
            .O(N__42453),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16 ));
    InMux I__9277 (
            .O(N__42450),
            .I(N__42446));
    InMux I__9276 (
            .O(N__42449),
            .I(N__42443));
    LocalMux I__9275 (
            .O(N__42446),
            .I(N__42439));
    LocalMux I__9274 (
            .O(N__42443),
            .I(N__42436));
    InMux I__9273 (
            .O(N__42442),
            .I(N__42433));
    Span12Mux_v I__9272 (
            .O(N__42439),
            .I(N__42430));
    Odrv4 I__9271 (
            .O(N__42436),
            .I(\delay_measurement_inst.N_363 ));
    LocalMux I__9270 (
            .O(N__42433),
            .I(\delay_measurement_inst.N_363 ));
    Odrv12 I__9269 (
            .O(N__42430),
            .I(\delay_measurement_inst.N_363 ));
    CascadeMux I__9268 (
            .O(N__42423),
            .I(N__42420));
    InMux I__9267 (
            .O(N__42420),
            .I(N__42417));
    LocalMux I__9266 (
            .O(N__42417),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0 ));
    CascadeMux I__9265 (
            .O(N__42414),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ));
    CascadeMux I__9264 (
            .O(N__42411),
            .I(elapsed_time_ns_1_RNIBA65M1_0_19_cascade_));
    CascadeMux I__9263 (
            .O(N__42408),
            .I(N__42405));
    InMux I__9262 (
            .O(N__42405),
            .I(N__42401));
    InMux I__9261 (
            .O(N__42404),
            .I(N__42398));
    LocalMux I__9260 (
            .O(N__42401),
            .I(N__42392));
    LocalMux I__9259 (
            .O(N__42398),
            .I(N__42392));
    InMux I__9258 (
            .O(N__42397),
            .I(N__42389));
    Span4Mux_h I__9257 (
            .O(N__42392),
            .I(N__42385));
    LocalMux I__9256 (
            .O(N__42389),
            .I(N__42382));
    InMux I__9255 (
            .O(N__42388),
            .I(N__42379));
    Odrv4 I__9254 (
            .O(N__42385),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ));
    Odrv4 I__9253 (
            .O(N__42382),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ));
    LocalMux I__9252 (
            .O(N__42379),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ));
    InMux I__9251 (
            .O(N__42372),
            .I(N__42369));
    LocalMux I__9250 (
            .O(N__42369),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20));
    CascadeMux I__9249 (
            .O(N__42366),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_));
    CascadeMux I__9248 (
            .O(N__42363),
            .I(N__42360));
    InMux I__9247 (
            .O(N__42360),
            .I(N__42357));
    LocalMux I__9246 (
            .O(N__42357),
            .I(N__42353));
    InMux I__9245 (
            .O(N__42356),
            .I(N__42350));
    Odrv4 I__9244 (
            .O(N__42353),
            .I(elapsed_time_ns_1_RNIRAIF91_0_21));
    LocalMux I__9243 (
            .O(N__42350),
            .I(elapsed_time_ns_1_RNIRAIF91_0_21));
    InMux I__9242 (
            .O(N__42345),
            .I(N__42342));
    LocalMux I__9241 (
            .O(N__42342),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15 ));
    CascadeMux I__9240 (
            .O(N__42339),
            .I(N__42336));
    InMux I__9239 (
            .O(N__42336),
            .I(N__42331));
    CascadeMux I__9238 (
            .O(N__42335),
            .I(N__42328));
    InMux I__9237 (
            .O(N__42334),
            .I(N__42325));
    LocalMux I__9236 (
            .O(N__42331),
            .I(N__42322));
    InMux I__9235 (
            .O(N__42328),
            .I(N__42318));
    LocalMux I__9234 (
            .O(N__42325),
            .I(N__42315));
    Span4Mux_h I__9233 (
            .O(N__42322),
            .I(N__42312));
    InMux I__9232 (
            .O(N__42321),
            .I(N__42309));
    LocalMux I__9231 (
            .O(N__42318),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    Odrv4 I__9230 (
            .O(N__42315),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    Odrv4 I__9229 (
            .O(N__42312),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    LocalMux I__9228 (
            .O(N__42309),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    InMux I__9227 (
            .O(N__42300),
            .I(N__42297));
    LocalMux I__9226 (
            .O(N__42297),
            .I(N__42294));
    Span4Mux_h I__9225 (
            .O(N__42294),
            .I(N__42291));
    Odrv4 I__9224 (
            .O(N__42291),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__9223 (
            .O(N__42288),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__9222 (
            .O(N__42285),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    CascadeMux I__9221 (
            .O(N__42282),
            .I(N__42279));
    InMux I__9220 (
            .O(N__42279),
            .I(N__42276));
    LocalMux I__9219 (
            .O(N__42276),
            .I(N__42273));
    Span4Mux_h I__9218 (
            .O(N__42273),
            .I(N__42270));
    Odrv4 I__9217 (
            .O(N__42270),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    CascadeMux I__9216 (
            .O(N__42267),
            .I(N__42263));
    CascadeMux I__9215 (
            .O(N__42266),
            .I(N__42260));
    InMux I__9214 (
            .O(N__42263),
            .I(N__42257));
    InMux I__9213 (
            .O(N__42260),
            .I(N__42254));
    LocalMux I__9212 (
            .O(N__42257),
            .I(N__42248));
    LocalMux I__9211 (
            .O(N__42254),
            .I(N__42248));
    CascadeMux I__9210 (
            .O(N__42253),
            .I(N__42245));
    Span4Mux_v I__9209 (
            .O(N__42248),
            .I(N__42242));
    InMux I__9208 (
            .O(N__42245),
            .I(N__42239));
    Odrv4 I__9207 (
            .O(N__42242),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    LocalMux I__9206 (
            .O(N__42239),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    InMux I__9205 (
            .O(N__42234),
            .I(N__42231));
    LocalMux I__9204 (
            .O(N__42231),
            .I(N__42226));
    InMux I__9203 (
            .O(N__42230),
            .I(N__42222));
    InMux I__9202 (
            .O(N__42229),
            .I(N__42219));
    Span12Mux_s11_v I__9201 (
            .O(N__42226),
            .I(N__42216));
    InMux I__9200 (
            .O(N__42225),
            .I(N__42213));
    LocalMux I__9199 (
            .O(N__42222),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__9198 (
            .O(N__42219),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    Odrv12 I__9197 (
            .O(N__42216),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__9196 (
            .O(N__42213),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    CascadeMux I__9195 (
            .O(N__42204),
            .I(N__42200));
    InMux I__9194 (
            .O(N__42203),
            .I(N__42196));
    InMux I__9193 (
            .O(N__42200),
            .I(N__42193));
    InMux I__9192 (
            .O(N__42199),
            .I(N__42190));
    LocalMux I__9191 (
            .O(N__42196),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    LocalMux I__9190 (
            .O(N__42193),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    LocalMux I__9189 (
            .O(N__42190),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    CascadeMux I__9188 (
            .O(N__42183),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10_cascade_));
    CascadeMux I__9187 (
            .O(N__42180),
            .I(N__42177));
    InMux I__9186 (
            .O(N__42177),
            .I(N__42174));
    LocalMux I__9185 (
            .O(N__42174),
            .I(N__42171));
    Span4Mux_v I__9184 (
            .O(N__42171),
            .I(N__42165));
    InMux I__9183 (
            .O(N__42170),
            .I(N__42162));
    InMux I__9182 (
            .O(N__42169),
            .I(N__42159));
    InMux I__9181 (
            .O(N__42168),
            .I(N__42155));
    Sp12to4 I__9180 (
            .O(N__42165),
            .I(N__42152));
    LocalMux I__9179 (
            .O(N__42162),
            .I(N__42149));
    LocalMux I__9178 (
            .O(N__42159),
            .I(N__42146));
    InMux I__9177 (
            .O(N__42158),
            .I(N__42143));
    LocalMux I__9176 (
            .O(N__42155),
            .I(elapsed_time_ns_1_RNI6565M1_0_14));
    Odrv12 I__9175 (
            .O(N__42152),
            .I(elapsed_time_ns_1_RNI6565M1_0_14));
    Odrv4 I__9174 (
            .O(N__42149),
            .I(elapsed_time_ns_1_RNI6565M1_0_14));
    Odrv4 I__9173 (
            .O(N__42146),
            .I(elapsed_time_ns_1_RNI6565M1_0_14));
    LocalMux I__9172 (
            .O(N__42143),
            .I(elapsed_time_ns_1_RNI6565M1_0_14));
    CascadeMux I__9171 (
            .O(N__42132),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_ ));
    InMux I__9170 (
            .O(N__42129),
            .I(N__42124));
    InMux I__9169 (
            .O(N__42128),
            .I(N__42120));
    InMux I__9168 (
            .O(N__42127),
            .I(N__42117));
    LocalMux I__9167 (
            .O(N__42124),
            .I(N__42114));
    InMux I__9166 (
            .O(N__42123),
            .I(N__42111));
    LocalMux I__9165 (
            .O(N__42120),
            .I(N__42106));
    LocalMux I__9164 (
            .O(N__42117),
            .I(N__42106));
    Span4Mux_v I__9163 (
            .O(N__42114),
            .I(N__42102));
    LocalMux I__9162 (
            .O(N__42111),
            .I(N__42097));
    Span4Mux_h I__9161 (
            .O(N__42106),
            .I(N__42097));
    InMux I__9160 (
            .O(N__42105),
            .I(N__42094));
    Odrv4 I__9159 (
            .O(N__42102),
            .I(elapsed_time_ns_1_RNIQENQL1_0_9));
    Odrv4 I__9158 (
            .O(N__42097),
            .I(elapsed_time_ns_1_RNIQENQL1_0_9));
    LocalMux I__9157 (
            .O(N__42094),
            .I(elapsed_time_ns_1_RNIQENQL1_0_9));
    CascadeMux I__9156 (
            .O(N__42087),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_ ));
    CascadeMux I__9155 (
            .O(N__42084),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ));
    CascadeMux I__9154 (
            .O(N__42081),
            .I(elapsed_time_ns_1_RNIK8NQL1_0_3_cascade_));
    CascadeMux I__9153 (
            .O(N__42078),
            .I(N__42075));
    InMux I__9152 (
            .O(N__42075),
            .I(N__42072));
    LocalMux I__9151 (
            .O(N__42072),
            .I(N__42069));
    Span4Mux_v I__9150 (
            .O(N__42069),
            .I(N__42066));
    Odrv4 I__9149 (
            .O(N__42066),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__9148 (
            .O(N__42063),
            .I(N__42060));
    LocalMux I__9147 (
            .O(N__42060),
            .I(N__42057));
    Span4Mux_h I__9146 (
            .O(N__42057),
            .I(N__42054));
    Odrv4 I__9145 (
            .O(N__42054),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__9144 (
            .O(N__42051),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__9143 (
            .O(N__42048),
            .I(N__42045));
    LocalMux I__9142 (
            .O(N__42045),
            .I(N__42042));
    Span4Mux_h I__9141 (
            .O(N__42042),
            .I(N__42039));
    Odrv4 I__9140 (
            .O(N__42039),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__9139 (
            .O(N__42036),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    CascadeMux I__9138 (
            .O(N__42033),
            .I(N__42030));
    InMux I__9137 (
            .O(N__42030),
            .I(N__42027));
    LocalMux I__9136 (
            .O(N__42027),
            .I(N__42024));
    Odrv12 I__9135 (
            .O(N__42024),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__9134 (
            .O(N__42021),
            .I(N__42018));
    LocalMux I__9133 (
            .O(N__42018),
            .I(N__42015));
    Span4Mux_h I__9132 (
            .O(N__42015),
            .I(N__42012));
    Odrv4 I__9131 (
            .O(N__42012),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__9130 (
            .O(N__42009),
            .I(bfn_17_14_0_));
    InMux I__9129 (
            .O(N__42006),
            .I(N__42003));
    LocalMux I__9128 (
            .O(N__42003),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__9127 (
            .O(N__42000),
            .I(N__41997));
    LocalMux I__9126 (
            .O(N__41997),
            .I(N__41994));
    Span4Mux_h I__9125 (
            .O(N__41994),
            .I(N__41991));
    Odrv4 I__9124 (
            .O(N__41991),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__9123 (
            .O(N__41988),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    CascadeMux I__9122 (
            .O(N__41985),
            .I(N__41982));
    InMux I__9121 (
            .O(N__41982),
            .I(N__41979));
    LocalMux I__9120 (
            .O(N__41979),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    CascadeMux I__9119 (
            .O(N__41976),
            .I(N__41973));
    InMux I__9118 (
            .O(N__41973),
            .I(N__41970));
    LocalMux I__9117 (
            .O(N__41970),
            .I(N__41967));
    Span4Mux_v I__9116 (
            .O(N__41967),
            .I(N__41964));
    Odrv4 I__9115 (
            .O(N__41964),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__9114 (
            .O(N__41961),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__9113 (
            .O(N__41958),
            .I(N__41955));
    LocalMux I__9112 (
            .O(N__41955),
            .I(N__41952));
    Span4Mux_v I__9111 (
            .O(N__41952),
            .I(N__41949));
    Odrv4 I__9110 (
            .O(N__41949),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__9109 (
            .O(N__41946),
            .I(N__41943));
    LocalMux I__9108 (
            .O(N__41943),
            .I(N__41940));
    Span4Mux_v I__9107 (
            .O(N__41940),
            .I(N__41937));
    Odrv4 I__9106 (
            .O(N__41937),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__9105 (
            .O(N__41934),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    CascadeMux I__9104 (
            .O(N__41931),
            .I(N__41928));
    InMux I__9103 (
            .O(N__41928),
            .I(N__41925));
    LocalMux I__9102 (
            .O(N__41925),
            .I(N__41922));
    Span4Mux_v I__9101 (
            .O(N__41922),
            .I(N__41919));
    Odrv4 I__9100 (
            .O(N__41919),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__9099 (
            .O(N__41916),
            .I(N__41913));
    LocalMux I__9098 (
            .O(N__41913),
            .I(N__41910));
    Span4Mux_h I__9097 (
            .O(N__41910),
            .I(N__41907));
    Odrv4 I__9096 (
            .O(N__41907),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__9095 (
            .O(N__41904),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__9094 (
            .O(N__41901),
            .I(N__41898));
    LocalMux I__9093 (
            .O(N__41898),
            .I(N__41895));
    Span4Mux_h I__9092 (
            .O(N__41895),
            .I(N__41892));
    Odrv4 I__9091 (
            .O(N__41892),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__9090 (
            .O(N__41889),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__9089 (
            .O(N__41886),
            .I(N__41883));
    LocalMux I__9088 (
            .O(N__41883),
            .I(N__41880));
    Span4Mux_v I__9087 (
            .O(N__41880),
            .I(N__41877));
    Odrv4 I__9086 (
            .O(N__41877),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__9085 (
            .O(N__41874),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__9084 (
            .O(N__41871),
            .I(N__41868));
    LocalMux I__9083 (
            .O(N__41868),
            .I(N__41865));
    Odrv4 I__9082 (
            .O(N__41865),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__9081 (
            .O(N__41862),
            .I(N__41859));
    LocalMux I__9080 (
            .O(N__41859),
            .I(N__41856));
    Span4Mux_h I__9079 (
            .O(N__41856),
            .I(N__41853));
    Odrv4 I__9078 (
            .O(N__41853),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__9077 (
            .O(N__41850),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__9076 (
            .O(N__41847),
            .I(N__41844));
    LocalMux I__9075 (
            .O(N__41844),
            .I(N__41841));
    Odrv12 I__9074 (
            .O(N__41841),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    InMux I__9073 (
            .O(N__41838),
            .I(N__41835));
    LocalMux I__9072 (
            .O(N__41835),
            .I(N__41832));
    Odrv12 I__9071 (
            .O(N__41832),
            .I(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ));
    InMux I__9070 (
            .O(N__41829),
            .I(N__41826));
    LocalMux I__9069 (
            .O(N__41826),
            .I(N__41823));
    Span4Mux_v I__9068 (
            .O(N__41823),
            .I(N__41820));
    Odrv4 I__9067 (
            .O(N__41820),
            .I(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ));
    InMux I__9066 (
            .O(N__41817),
            .I(N__41814));
    LocalMux I__9065 (
            .O(N__41814),
            .I(N__41811));
    Odrv4 I__9064 (
            .O(N__41811),
            .I(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ));
    CascadeMux I__9063 (
            .O(N__41808),
            .I(N__41805));
    InMux I__9062 (
            .O(N__41805),
            .I(N__41802));
    LocalMux I__9061 (
            .O(N__41802),
            .I(N__41799));
    Odrv12 I__9060 (
            .O(N__41799),
            .I(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ));
    InMux I__9059 (
            .O(N__41796),
            .I(N__41793));
    LocalMux I__9058 (
            .O(N__41793),
            .I(N__41790));
    Odrv12 I__9057 (
            .O(N__41790),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__9056 (
            .O(N__41787),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__9055 (
            .O(N__41784),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__9054 (
            .O(N__41781),
            .I(N__41777));
    CascadeMux I__9053 (
            .O(N__41780),
            .I(N__41774));
    InMux I__9052 (
            .O(N__41777),
            .I(N__41771));
    InMux I__9051 (
            .O(N__41774),
            .I(N__41768));
    LocalMux I__9050 (
            .O(N__41771),
            .I(N__41765));
    LocalMux I__9049 (
            .O(N__41768),
            .I(N__41762));
    Span4Mux_v I__9048 (
            .O(N__41765),
            .I(N__41756));
    Span4Mux_h I__9047 (
            .O(N__41762),
            .I(N__41756));
    CascadeMux I__9046 (
            .O(N__41761),
            .I(N__41753));
    Span4Mux_h I__9045 (
            .O(N__41756),
            .I(N__41749));
    InMux I__9044 (
            .O(N__41753),
            .I(N__41744));
    InMux I__9043 (
            .O(N__41752),
            .I(N__41744));
    Odrv4 I__9042 (
            .O(N__41749),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__9041 (
            .O(N__41744),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__9040 (
            .O(N__41739),
            .I(N__41736));
    LocalMux I__9039 (
            .O(N__41736),
            .I(N__41731));
    InMux I__9038 (
            .O(N__41735),
            .I(N__41728));
    InMux I__9037 (
            .O(N__41734),
            .I(N__41725));
    Span4Mux_v I__9036 (
            .O(N__41731),
            .I(N__41720));
    LocalMux I__9035 (
            .O(N__41728),
            .I(N__41720));
    LocalMux I__9034 (
            .O(N__41725),
            .I(N__41717));
    Span4Mux_h I__9033 (
            .O(N__41720),
            .I(N__41714));
    Odrv4 I__9032 (
            .O(N__41717),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__9031 (
            .O(N__41714),
            .I(\current_shift_inst.un4_control_input1_12 ));
    CascadeMux I__9030 (
            .O(N__41709),
            .I(N__41705));
    InMux I__9029 (
            .O(N__41708),
            .I(N__41702));
    InMux I__9028 (
            .O(N__41705),
            .I(N__41698));
    LocalMux I__9027 (
            .O(N__41702),
            .I(N__41694));
    InMux I__9026 (
            .O(N__41701),
            .I(N__41691));
    LocalMux I__9025 (
            .O(N__41698),
            .I(N__41688));
    InMux I__9024 (
            .O(N__41697),
            .I(N__41685));
    Span4Mux_v I__9023 (
            .O(N__41694),
            .I(N__41680));
    LocalMux I__9022 (
            .O(N__41691),
            .I(N__41680));
    Span4Mux_v I__9021 (
            .O(N__41688),
            .I(N__41677));
    LocalMux I__9020 (
            .O(N__41685),
            .I(N__41674));
    Span4Mux_h I__9019 (
            .O(N__41680),
            .I(N__41671));
    Span4Mux_h I__9018 (
            .O(N__41677),
            .I(N__41666));
    Span4Mux_h I__9017 (
            .O(N__41674),
            .I(N__41666));
    Odrv4 I__9016 (
            .O(N__41671),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__9015 (
            .O(N__41666),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__9014 (
            .O(N__41661),
            .I(N__41658));
    LocalMux I__9013 (
            .O(N__41658),
            .I(N__41653));
    InMux I__9012 (
            .O(N__41657),
            .I(N__41650));
    InMux I__9011 (
            .O(N__41656),
            .I(N__41647));
    Span4Mux_v I__9010 (
            .O(N__41653),
            .I(N__41642));
    LocalMux I__9009 (
            .O(N__41650),
            .I(N__41642));
    LocalMux I__9008 (
            .O(N__41647),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv4 I__9007 (
            .O(N__41642),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__9006 (
            .O(N__41637),
            .I(N__41634));
    LocalMux I__9005 (
            .O(N__41634),
            .I(N__41630));
    InMux I__9004 (
            .O(N__41633),
            .I(N__41627));
    Span4Mux_h I__9003 (
            .O(N__41630),
            .I(N__41624));
    LocalMux I__9002 (
            .O(N__41627),
            .I(N__41621));
    Odrv4 I__9001 (
            .O(N__41624),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    Odrv4 I__9000 (
            .O(N__41621),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    InMux I__8999 (
            .O(N__41616),
            .I(N__41613));
    LocalMux I__8998 (
            .O(N__41613),
            .I(N__41609));
    CascadeMux I__8997 (
            .O(N__41612),
            .I(N__41606));
    Span4Mux_v I__8996 (
            .O(N__41609),
            .I(N__41603));
    InMux I__8995 (
            .O(N__41606),
            .I(N__41600));
    Odrv4 I__8994 (
            .O(N__41603),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    LocalMux I__8993 (
            .O(N__41600),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__8992 (
            .O(N__41595),
            .I(N__41592));
    InMux I__8991 (
            .O(N__41592),
            .I(N__41589));
    LocalMux I__8990 (
            .O(N__41589),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__8989 (
            .O(N__41586),
            .I(N__41583));
    LocalMux I__8988 (
            .O(N__41583),
            .I(N__41580));
    Span4Mux_v I__8987 (
            .O(N__41580),
            .I(N__41577));
    Odrv4 I__8986 (
            .O(N__41577),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    CascadeMux I__8985 (
            .O(N__41574),
            .I(N__41571));
    InMux I__8984 (
            .O(N__41571),
            .I(N__41568));
    LocalMux I__8983 (
            .O(N__41568),
            .I(N__41565));
    Span4Mux_v I__8982 (
            .O(N__41565),
            .I(N__41562));
    Odrv4 I__8981 (
            .O(N__41562),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    InMux I__8980 (
            .O(N__41559),
            .I(N__41556));
    LocalMux I__8979 (
            .O(N__41556),
            .I(N__41553));
    Odrv4 I__8978 (
            .O(N__41553),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__8977 (
            .O(N__41550),
            .I(N__41541));
    InMux I__8976 (
            .O(N__41549),
            .I(N__41541));
    InMux I__8975 (
            .O(N__41548),
            .I(N__41541));
    LocalMux I__8974 (
            .O(N__41541),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__8973 (
            .O(N__41538),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__8972 (
            .O(N__41535),
            .I(N__41532));
    LocalMux I__8971 (
            .O(N__41532),
            .I(N__41529));
    Odrv4 I__8970 (
            .O(N__41529),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__8969 (
            .O(N__41526),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__8968 (
            .O(N__41523),
            .I(N__41520));
    LocalMux I__8967 (
            .O(N__41520),
            .I(N__41517));
    Odrv4 I__8966 (
            .O(N__41517),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__8965 (
            .O(N__41514),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__8964 (
            .O(N__41511),
            .I(N__41508));
    LocalMux I__8963 (
            .O(N__41508),
            .I(N__41505));
    Span4Mux_h I__8962 (
            .O(N__41505),
            .I(N__41502));
    Span4Mux_h I__8961 (
            .O(N__41502),
            .I(N__41499));
    Odrv4 I__8960 (
            .O(N__41499),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__8959 (
            .O(N__41496),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__8958 (
            .O(N__41493),
            .I(N__41490));
    LocalMux I__8957 (
            .O(N__41490),
            .I(N__41487));
    Odrv4 I__8956 (
            .O(N__41487),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    CascadeMux I__8955 (
            .O(N__41484),
            .I(N__41481));
    InMux I__8954 (
            .O(N__41481),
            .I(N__41477));
    InMux I__8953 (
            .O(N__41480),
            .I(N__41474));
    LocalMux I__8952 (
            .O(N__41477),
            .I(N__41468));
    LocalMux I__8951 (
            .O(N__41474),
            .I(N__41468));
    InMux I__8950 (
            .O(N__41473),
            .I(N__41465));
    Span4Mux_v I__8949 (
            .O(N__41468),
            .I(N__41462));
    LocalMux I__8948 (
            .O(N__41465),
            .I(N__41459));
    Odrv4 I__8947 (
            .O(N__41462),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv12 I__8946 (
            .O(N__41459),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__8945 (
            .O(N__41454),
            .I(bfn_17_10_0_));
    InMux I__8944 (
            .O(N__41451),
            .I(N__41448));
    LocalMux I__8943 (
            .O(N__41448),
            .I(N__41445));
    Odrv12 I__8942 (
            .O(N__41445),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    CascadeMux I__8941 (
            .O(N__41442),
            .I(N__41439));
    InMux I__8940 (
            .O(N__41439),
            .I(N__41435));
    InMux I__8939 (
            .O(N__41438),
            .I(N__41432));
    LocalMux I__8938 (
            .O(N__41435),
            .I(N__41428));
    LocalMux I__8937 (
            .O(N__41432),
            .I(N__41425));
    InMux I__8936 (
            .O(N__41431),
            .I(N__41422));
    Sp12to4 I__8935 (
            .O(N__41428),
            .I(N__41419));
    Span4Mux_v I__8934 (
            .O(N__41425),
            .I(N__41414));
    LocalMux I__8933 (
            .O(N__41422),
            .I(N__41414));
    Odrv12 I__8932 (
            .O(N__41419),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__8931 (
            .O(N__41414),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__8930 (
            .O(N__41409),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__8929 (
            .O(N__41406),
            .I(N__41403));
    LocalMux I__8928 (
            .O(N__41403),
            .I(N__41400));
    Odrv12 I__8927 (
            .O(N__41400),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    CascadeMux I__8926 (
            .O(N__41397),
            .I(N__41394));
    InMux I__8925 (
            .O(N__41394),
            .I(N__41391));
    LocalMux I__8924 (
            .O(N__41391),
            .I(N__41387));
    CascadeMux I__8923 (
            .O(N__41390),
            .I(N__41384));
    Span4Mux_v I__8922 (
            .O(N__41387),
            .I(N__41380));
    InMux I__8921 (
            .O(N__41384),
            .I(N__41375));
    InMux I__8920 (
            .O(N__41383),
            .I(N__41375));
    Odrv4 I__8919 (
            .O(N__41380),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__8918 (
            .O(N__41375),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__8917 (
            .O(N__41370),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__8916 (
            .O(N__41367),
            .I(N__41364));
    LocalMux I__8915 (
            .O(N__41364),
            .I(N__41361));
    Odrv12 I__8914 (
            .O(N__41361),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__8913 (
            .O(N__41358),
            .I(N__41349));
    InMux I__8912 (
            .O(N__41357),
            .I(N__41349));
    InMux I__8911 (
            .O(N__41356),
            .I(N__41349));
    LocalMux I__8910 (
            .O(N__41349),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__8909 (
            .O(N__41346),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__8908 (
            .O(N__41343),
            .I(N__41340));
    LocalMux I__8907 (
            .O(N__41340),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__8906 (
            .O(N__41337),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__8905 (
            .O(N__41334),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__8904 (
            .O(N__41331),
            .I(N__41328));
    LocalMux I__8903 (
            .O(N__41328),
            .I(N__41325));
    Span4Mux_h I__8902 (
            .O(N__41325),
            .I(N__41322));
    Odrv4 I__8901 (
            .O(N__41322),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__8900 (
            .O(N__41319),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__8899 (
            .O(N__41316),
            .I(N__41313));
    LocalMux I__8898 (
            .O(N__41313),
            .I(N__41310));
    Odrv12 I__8897 (
            .O(N__41310),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__8896 (
            .O(N__41307),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__8895 (
            .O(N__41304),
            .I(N__41301));
    LocalMux I__8894 (
            .O(N__41301),
            .I(N__41298));
    Odrv4 I__8893 (
            .O(N__41298),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__8892 (
            .O(N__41295),
            .I(bfn_17_9_0_));
    InMux I__8891 (
            .O(N__41292),
            .I(N__41289));
    LocalMux I__8890 (
            .O(N__41289),
            .I(N__41286));
    Odrv12 I__8889 (
            .O(N__41286),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__8888 (
            .O(N__41283),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__8887 (
            .O(N__41280),
            .I(N__41277));
    LocalMux I__8886 (
            .O(N__41277),
            .I(N__41274));
    Odrv12 I__8885 (
            .O(N__41274),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__8884 (
            .O(N__41271),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__8883 (
            .O(N__41268),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__8882 (
            .O(N__41265),
            .I(N__41262));
    LocalMux I__8881 (
            .O(N__41262),
            .I(N__41259));
    Odrv4 I__8880 (
            .O(N__41259),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__8879 (
            .O(N__41256),
            .I(N__41253));
    LocalMux I__8878 (
            .O(N__41253),
            .I(N__41248));
    InMux I__8877 (
            .O(N__41252),
            .I(N__41245));
    InMux I__8876 (
            .O(N__41251),
            .I(N__41242));
    Odrv4 I__8875 (
            .O(N__41248),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__8874 (
            .O(N__41245),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__8873 (
            .O(N__41242),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__8872 (
            .O(N__41235),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__8871 (
            .O(N__41232),
            .I(N__41229));
    LocalMux I__8870 (
            .O(N__41229),
            .I(N__41226));
    Span4Mux_h I__8869 (
            .O(N__41226),
            .I(N__41223));
    Odrv4 I__8868 (
            .O(N__41223),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__8867 (
            .O(N__41220),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__8866 (
            .O(N__41217),
            .I(N__41214));
    LocalMux I__8865 (
            .O(N__41214),
            .I(N__41211));
    Odrv4 I__8864 (
            .O(N__41211),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__8863 (
            .O(N__41208),
            .I(N__41205));
    LocalMux I__8862 (
            .O(N__41205),
            .I(N__41200));
    InMux I__8861 (
            .O(N__41204),
            .I(N__41197));
    InMux I__8860 (
            .O(N__41203),
            .I(N__41194));
    Span4Mux_v I__8859 (
            .O(N__41200),
            .I(N__41189));
    LocalMux I__8858 (
            .O(N__41197),
            .I(N__41189));
    LocalMux I__8857 (
            .O(N__41194),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__8856 (
            .O(N__41189),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__8855 (
            .O(N__41184),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__8854 (
            .O(N__41181),
            .I(N__41178));
    LocalMux I__8853 (
            .O(N__41178),
            .I(N__41175));
    Odrv4 I__8852 (
            .O(N__41175),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__8851 (
            .O(N__41172),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__8850 (
            .O(N__41169),
            .I(N__41166));
    LocalMux I__8849 (
            .O(N__41166),
            .I(N__41163));
    Span4Mux_h I__8848 (
            .O(N__41163),
            .I(N__41160));
    Odrv4 I__8847 (
            .O(N__41160),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__8846 (
            .O(N__41157),
            .I(N__41153));
    CascadeMux I__8845 (
            .O(N__41156),
            .I(N__41150));
    LocalMux I__8844 (
            .O(N__41153),
            .I(N__41146));
    InMux I__8843 (
            .O(N__41150),
            .I(N__41141));
    InMux I__8842 (
            .O(N__41149),
            .I(N__41141));
    Span4Mux_h I__8841 (
            .O(N__41146),
            .I(N__41138));
    LocalMux I__8840 (
            .O(N__41141),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv4 I__8839 (
            .O(N__41138),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__8838 (
            .O(N__41133),
            .I(bfn_17_8_0_));
    InMux I__8837 (
            .O(N__41130),
            .I(N__41127));
    LocalMux I__8836 (
            .O(N__41127),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__8835 (
            .O(N__41124),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__8834 (
            .O(N__41121),
            .I(N__41118));
    LocalMux I__8833 (
            .O(N__41118),
            .I(N__41115));
    Span4Mux_h I__8832 (
            .O(N__41115),
            .I(N__41112));
    Odrv4 I__8831 (
            .O(N__41112),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__8830 (
            .O(N__41109),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__8829 (
            .O(N__41106),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    CascadeMux I__8828 (
            .O(N__41103),
            .I(N__41099));
    CascadeMux I__8827 (
            .O(N__41102),
            .I(N__41096));
    InMux I__8826 (
            .O(N__41099),
            .I(N__41093));
    InMux I__8825 (
            .O(N__41096),
            .I(N__41090));
    LocalMux I__8824 (
            .O(N__41093),
            .I(N__41085));
    LocalMux I__8823 (
            .O(N__41090),
            .I(N__41082));
    InMux I__8822 (
            .O(N__41089),
            .I(N__41077));
    InMux I__8821 (
            .O(N__41088),
            .I(N__41077));
    Span4Mux_h I__8820 (
            .O(N__41085),
            .I(N__41074));
    Span4Mux_v I__8819 (
            .O(N__41082),
            .I(N__41069));
    LocalMux I__8818 (
            .O(N__41077),
            .I(N__41069));
    Odrv4 I__8817 (
            .O(N__41074),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__8816 (
            .O(N__41069),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__8815 (
            .O(N__41064),
            .I(N__41060));
    InMux I__8814 (
            .O(N__41063),
            .I(N__41057));
    LocalMux I__8813 (
            .O(N__41060),
            .I(N__41053));
    LocalMux I__8812 (
            .O(N__41057),
            .I(N__41050));
    CascadeMux I__8811 (
            .O(N__41056),
            .I(N__41046));
    Span4Mux_h I__8810 (
            .O(N__41053),
            .I(N__41041));
    Span4Mux_v I__8809 (
            .O(N__41050),
            .I(N__41041));
    InMux I__8808 (
            .O(N__41049),
            .I(N__41038));
    InMux I__8807 (
            .O(N__41046),
            .I(N__41035));
    Odrv4 I__8806 (
            .O(N__41041),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__8805 (
            .O(N__41038),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__8804 (
            .O(N__41035),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__8803 (
            .O(N__41028),
            .I(N__41025));
    LocalMux I__8802 (
            .O(N__41025),
            .I(N__41022));
    Odrv4 I__8801 (
            .O(N__41022),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__8800 (
            .O(N__41019),
            .I(N__41013));
    InMux I__8799 (
            .O(N__41018),
            .I(N__41013));
    LocalMux I__8798 (
            .O(N__41013),
            .I(N__41010));
    Span4Mux_v I__8797 (
            .O(N__41010),
            .I(N__41006));
    InMux I__8796 (
            .O(N__41009),
            .I(N__41003));
    Odrv4 I__8795 (
            .O(N__41006),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__8794 (
            .O(N__41003),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__8793 (
            .O(N__40998),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__8792 (
            .O(N__40995),
            .I(N__40992));
    LocalMux I__8791 (
            .O(N__40992),
            .I(N__40989));
    Odrv12 I__8790 (
            .O(N__40989),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__8789 (
            .O(N__40986),
            .I(N__40983));
    LocalMux I__8788 (
            .O(N__40983),
            .I(N__40980));
    Span4Mux_v I__8787 (
            .O(N__40980),
            .I(N__40975));
    InMux I__8786 (
            .O(N__40979),
            .I(N__40972));
    InMux I__8785 (
            .O(N__40978),
            .I(N__40969));
    Odrv4 I__8784 (
            .O(N__40975),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__8783 (
            .O(N__40972),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__8782 (
            .O(N__40969),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__8781 (
            .O(N__40962),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__8780 (
            .O(N__40959),
            .I(N__40956));
    LocalMux I__8779 (
            .O(N__40956),
            .I(N__40953));
    Odrv4 I__8778 (
            .O(N__40953),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    CascadeMux I__8777 (
            .O(N__40950),
            .I(N__40947));
    InMux I__8776 (
            .O(N__40947),
            .I(N__40944));
    LocalMux I__8775 (
            .O(N__40944),
            .I(N__40939));
    InMux I__8774 (
            .O(N__40943),
            .I(N__40934));
    InMux I__8773 (
            .O(N__40942),
            .I(N__40934));
    Span4Mux_h I__8772 (
            .O(N__40939),
            .I(N__40931));
    LocalMux I__8771 (
            .O(N__40934),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__8770 (
            .O(N__40931),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__8769 (
            .O(N__40926),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__8768 (
            .O(N__40923),
            .I(N__40918));
    InMux I__8767 (
            .O(N__40922),
            .I(N__40915));
    InMux I__8766 (
            .O(N__40921),
            .I(N__40911));
    LocalMux I__8765 (
            .O(N__40918),
            .I(N__40908));
    LocalMux I__8764 (
            .O(N__40915),
            .I(N__40905));
    InMux I__8763 (
            .O(N__40914),
            .I(N__40902));
    LocalMux I__8762 (
            .O(N__40911),
            .I(N__40899));
    Span12Mux_v I__8761 (
            .O(N__40908),
            .I(N__40896));
    Span12Mux_v I__8760 (
            .O(N__40905),
            .I(N__40893));
    LocalMux I__8759 (
            .O(N__40902),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__8758 (
            .O(N__40899),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv12 I__8757 (
            .O(N__40896),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv12 I__8756 (
            .O(N__40893),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__8755 (
            .O(N__40884),
            .I(N__40881));
    LocalMux I__8754 (
            .O(N__40881),
            .I(N__40878));
    Span4Mux_h I__8753 (
            .O(N__40878),
            .I(N__40875));
    Odrv4 I__8752 (
            .O(N__40875),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5 ));
    CascadeMux I__8751 (
            .O(N__40872),
            .I(N__40869));
    InMux I__8750 (
            .O(N__40869),
            .I(N__40861));
    InMux I__8749 (
            .O(N__40868),
            .I(N__40855));
    InMux I__8748 (
            .O(N__40867),
            .I(N__40850));
    InMux I__8747 (
            .O(N__40866),
            .I(N__40850));
    InMux I__8746 (
            .O(N__40865),
            .I(N__40845));
    InMux I__8745 (
            .O(N__40864),
            .I(N__40845));
    LocalMux I__8744 (
            .O(N__40861),
            .I(N__40842));
    CascadeMux I__8743 (
            .O(N__40860),
            .I(N__40839));
    CascadeMux I__8742 (
            .O(N__40859),
            .I(N__40835));
    CascadeMux I__8741 (
            .O(N__40858),
            .I(N__40832));
    LocalMux I__8740 (
            .O(N__40855),
            .I(N__40828));
    LocalMux I__8739 (
            .O(N__40850),
            .I(N__40825));
    LocalMux I__8738 (
            .O(N__40845),
            .I(N__40820));
    Span4Mux_v I__8737 (
            .O(N__40842),
            .I(N__40820));
    InMux I__8736 (
            .O(N__40839),
            .I(N__40815));
    InMux I__8735 (
            .O(N__40838),
            .I(N__40815));
    InMux I__8734 (
            .O(N__40835),
            .I(N__40812));
    InMux I__8733 (
            .O(N__40832),
            .I(N__40807));
    InMux I__8732 (
            .O(N__40831),
            .I(N__40807));
    Span4Mux_h I__8731 (
            .O(N__40828),
            .I(N__40804));
    Span4Mux_v I__8730 (
            .O(N__40825),
            .I(N__40801));
    Span4Mux_v I__8729 (
            .O(N__40820),
            .I(N__40798));
    LocalMux I__8728 (
            .O(N__40815),
            .I(\phase_controller_inst1.stoper_tr.N_242 ));
    LocalMux I__8727 (
            .O(N__40812),
            .I(\phase_controller_inst1.stoper_tr.N_242 ));
    LocalMux I__8726 (
            .O(N__40807),
            .I(\phase_controller_inst1.stoper_tr.N_242 ));
    Odrv4 I__8725 (
            .O(N__40804),
            .I(\phase_controller_inst1.stoper_tr.N_242 ));
    Odrv4 I__8724 (
            .O(N__40801),
            .I(\phase_controller_inst1.stoper_tr.N_242 ));
    Odrv4 I__8723 (
            .O(N__40798),
            .I(\phase_controller_inst1.stoper_tr.N_242 ));
    InMux I__8722 (
            .O(N__40785),
            .I(N__40782));
    LocalMux I__8721 (
            .O(N__40782),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__8720 (
            .O(N__40779),
            .I(N__40776));
    InMux I__8719 (
            .O(N__40776),
            .I(N__40770));
    InMux I__8718 (
            .O(N__40775),
            .I(N__40770));
    LocalMux I__8717 (
            .O(N__40770),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__8716 (
            .O(N__40767),
            .I(N__40763));
    CascadeMux I__8715 (
            .O(N__40766),
            .I(N__40760));
    InMux I__8714 (
            .O(N__40763),
            .I(N__40757));
    InMux I__8713 (
            .O(N__40760),
            .I(N__40754));
    LocalMux I__8712 (
            .O(N__40757),
            .I(N__40751));
    LocalMux I__8711 (
            .O(N__40754),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    Odrv4 I__8710 (
            .O(N__40751),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__8709 (
            .O(N__40746),
            .I(N__40742));
    InMux I__8708 (
            .O(N__40745),
            .I(N__40739));
    LocalMux I__8707 (
            .O(N__40742),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    LocalMux I__8706 (
            .O(N__40739),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__8705 (
            .O(N__40734),
            .I(N__40730));
    InMux I__8704 (
            .O(N__40733),
            .I(N__40727));
    LocalMux I__8703 (
            .O(N__40730),
            .I(N__40723));
    LocalMux I__8702 (
            .O(N__40727),
            .I(N__40720));
    InMux I__8701 (
            .O(N__40726),
            .I(N__40717));
    Span4Mux_h I__8700 (
            .O(N__40723),
            .I(N__40714));
    Odrv4 I__8699 (
            .O(N__40720),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__8698 (
            .O(N__40717),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__8697 (
            .O(N__40714),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    CascadeMux I__8696 (
            .O(N__40707),
            .I(N__40704));
    InMux I__8695 (
            .O(N__40704),
            .I(N__40699));
    InMux I__8694 (
            .O(N__40703),
            .I(N__40696));
    CascadeMux I__8693 (
            .O(N__40702),
            .I(N__40693));
    LocalMux I__8692 (
            .O(N__40699),
            .I(N__40689));
    LocalMux I__8691 (
            .O(N__40696),
            .I(N__40686));
    InMux I__8690 (
            .O(N__40693),
            .I(N__40681));
    InMux I__8689 (
            .O(N__40692),
            .I(N__40681));
    Span4Mux_v I__8688 (
            .O(N__40689),
            .I(N__40678));
    Span4Mux_h I__8687 (
            .O(N__40686),
            .I(N__40673));
    LocalMux I__8686 (
            .O(N__40681),
            .I(N__40673));
    Odrv4 I__8685 (
            .O(N__40678),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__8684 (
            .O(N__40673),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__8683 (
            .O(N__40668),
            .I(N__40661));
    InMux I__8682 (
            .O(N__40667),
            .I(N__40661));
    InMux I__8681 (
            .O(N__40666),
            .I(N__40658));
    LocalMux I__8680 (
            .O(N__40661),
            .I(N__40655));
    LocalMux I__8679 (
            .O(N__40658),
            .I(N__40652));
    Span4Mux_v I__8678 (
            .O(N__40655),
            .I(N__40648));
    Span4Mux_v I__8677 (
            .O(N__40652),
            .I(N__40645));
    InMux I__8676 (
            .O(N__40651),
            .I(N__40642));
    Odrv4 I__8675 (
            .O(N__40648),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    Odrv4 I__8674 (
            .O(N__40645),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__8673 (
            .O(N__40642),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__8672 (
            .O(N__40635),
            .I(N__40632));
    InMux I__8671 (
            .O(N__40632),
            .I(N__40628));
    InMux I__8670 (
            .O(N__40631),
            .I(N__40625));
    LocalMux I__8669 (
            .O(N__40628),
            .I(\delay_measurement_inst.delay_tr_timer.N_382 ));
    LocalMux I__8668 (
            .O(N__40625),
            .I(\delay_measurement_inst.delay_tr_timer.N_382 ));
    CascadeMux I__8667 (
            .O(N__40620),
            .I(\delay_measurement_inst.delay_tr_timer.N_382_cascade_ ));
    InMux I__8666 (
            .O(N__40617),
            .I(N__40613));
    InMux I__8665 (
            .O(N__40616),
            .I(N__40610));
    LocalMux I__8664 (
            .O(N__40613),
            .I(\delay_measurement_inst.delay_tr_timer.N_371 ));
    LocalMux I__8663 (
            .O(N__40610),
            .I(\delay_measurement_inst.delay_tr_timer.N_371 ));
    InMux I__8662 (
            .O(N__40605),
            .I(N__40599));
    InMux I__8661 (
            .O(N__40604),
            .I(N__40599));
    LocalMux I__8660 (
            .O(N__40599),
            .I(\delay_measurement_inst.delay_tr_timer.N_356 ));
    InMux I__8659 (
            .O(N__40596),
            .I(N__40593));
    LocalMux I__8658 (
            .O(N__40593),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ));
    CascadeMux I__8657 (
            .O(N__40590),
            .I(\delay_measurement_inst.delay_tr_timer.N_351_cascade_ ));
    InMux I__8656 (
            .O(N__40587),
            .I(N__40583));
    CascadeMux I__8655 (
            .O(N__40586),
            .I(N__40580));
    LocalMux I__8654 (
            .O(N__40583),
            .I(N__40577));
    InMux I__8653 (
            .O(N__40580),
            .I(N__40574));
    Odrv4 I__8652 (
            .O(N__40577),
            .I(\delay_measurement_inst.delay_tr_timer.N_378 ));
    LocalMux I__8651 (
            .O(N__40574),
            .I(\delay_measurement_inst.delay_tr_timer.N_378 ));
    InMux I__8650 (
            .O(N__40569),
            .I(N__40566));
    LocalMux I__8649 (
            .O(N__40566),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4 ));
    InMux I__8648 (
            .O(N__40563),
            .I(N__40560));
    LocalMux I__8647 (
            .O(N__40560),
            .I(N__40556));
    InMux I__8646 (
            .O(N__40559),
            .I(N__40553));
    Odrv4 I__8645 (
            .O(N__40556),
            .I(\delay_measurement_inst.delay_tr_timer.N_360 ));
    LocalMux I__8644 (
            .O(N__40553),
            .I(\delay_measurement_inst.delay_tr_timer.N_360 ));
    CascadeMux I__8643 (
            .O(N__40548),
            .I(\delay_measurement_inst.delay_tr9_cascade_ ));
    InMux I__8642 (
            .O(N__40545),
            .I(N__40542));
    LocalMux I__8641 (
            .O(N__40542),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0 ));
    InMux I__8640 (
            .O(N__40539),
            .I(N__40533));
    InMux I__8639 (
            .O(N__40538),
            .I(N__40533));
    LocalMux I__8638 (
            .O(N__40533),
            .I(\delay_measurement_inst.delay_tr_timer.N_390 ));
    CascadeMux I__8637 (
            .O(N__40530),
            .I(\delay_measurement_inst.delay_tr_timer.N_390_cascade_ ));
    CascadeMux I__8636 (
            .O(N__40527),
            .I(\delay_measurement_inst.delay_tr_timer.N_391_cascade_ ));
    CascadeMux I__8635 (
            .O(N__40524),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ));
    CascadeMux I__8634 (
            .O(N__40521),
            .I(elapsed_time_ns_1_RNI6565M1_0_14_cascade_));
    InMux I__8633 (
            .O(N__40518),
            .I(N__40515));
    LocalMux I__8632 (
            .O(N__40515),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14 ));
    InMux I__8631 (
            .O(N__40512),
            .I(N__40509));
    LocalMux I__8630 (
            .O(N__40509),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25));
    InMux I__8629 (
            .O(N__40506),
            .I(N__40500));
    InMux I__8628 (
            .O(N__40505),
            .I(N__40500));
    LocalMux I__8627 (
            .O(N__40500),
            .I(elapsed_time_ns_1_RNI1HIF91_0_27));
    CascadeMux I__8626 (
            .O(N__40497),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_));
    InMux I__8625 (
            .O(N__40494),
            .I(N__40488));
    InMux I__8624 (
            .O(N__40493),
            .I(N__40488));
    LocalMux I__8623 (
            .O(N__40488),
            .I(elapsed_time_ns_1_RNISBIF91_0_22));
    CascadeMux I__8622 (
            .O(N__40485),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15_cascade_ ));
    InMux I__8621 (
            .O(N__40482),
            .I(N__40476));
    InMux I__8620 (
            .O(N__40481),
            .I(N__40476));
    LocalMux I__8619 (
            .O(N__40476),
            .I(elapsed_time_ns_1_RNI2IIF91_0_28));
    CascadeMux I__8618 (
            .O(N__40473),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ));
    InMux I__8617 (
            .O(N__40470),
            .I(N__40466));
    InMux I__8616 (
            .O(N__40469),
            .I(N__40463));
    LocalMux I__8615 (
            .O(N__40466),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    LocalMux I__8614 (
            .O(N__40463),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    InMux I__8613 (
            .O(N__40458),
            .I(N__40455));
    LocalMux I__8612 (
            .O(N__40455),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ));
    InMux I__8611 (
            .O(N__40452),
            .I(N__40449));
    LocalMux I__8610 (
            .O(N__40449),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ));
    InMux I__8609 (
            .O(N__40446),
            .I(N__40442));
    InMux I__8608 (
            .O(N__40445),
            .I(N__40439));
    LocalMux I__8607 (
            .O(N__40442),
            .I(N__40434));
    LocalMux I__8606 (
            .O(N__40439),
            .I(N__40434));
    Span4Mux_h I__8605 (
            .O(N__40434),
            .I(N__40430));
    InMux I__8604 (
            .O(N__40433),
            .I(N__40427));
    Span4Mux_h I__8603 (
            .O(N__40430),
            .I(N__40424));
    LocalMux I__8602 (
            .O(N__40427),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    Odrv4 I__8601 (
            .O(N__40424),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    InMux I__8600 (
            .O(N__40419),
            .I(N__40416));
    LocalMux I__8599 (
            .O(N__40416),
            .I(N__40411));
    InMux I__8598 (
            .O(N__40415),
            .I(N__40408));
    InMux I__8597 (
            .O(N__40414),
            .I(N__40405));
    Span4Mux_v I__8596 (
            .O(N__40411),
            .I(N__40398));
    LocalMux I__8595 (
            .O(N__40408),
            .I(N__40398));
    LocalMux I__8594 (
            .O(N__40405),
            .I(N__40398));
    Span4Mux_h I__8593 (
            .O(N__40398),
            .I(N__40394));
    InMux I__8592 (
            .O(N__40397),
            .I(N__40391));
    Odrv4 I__8591 (
            .O(N__40394),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__8590 (
            .O(N__40391),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__8589 (
            .O(N__40386),
            .I(N__40383));
    LocalMux I__8588 (
            .O(N__40383),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    CascadeMux I__8587 (
            .O(N__40380),
            .I(elapsed_time_ns_1_RNISAHF91_0_13_cascade_));
    InMux I__8586 (
            .O(N__40377),
            .I(N__40374));
    LocalMux I__8585 (
            .O(N__40374),
            .I(N__40371));
    Span4Mux_v I__8584 (
            .O(N__40371),
            .I(N__40368));
    Odrv4 I__8583 (
            .O(N__40368),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__8582 (
            .O(N__40365),
            .I(N__40362));
    LocalMux I__8581 (
            .O(N__40362),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ));
    InMux I__8580 (
            .O(N__40359),
            .I(N__40356));
    LocalMux I__8579 (
            .O(N__40356),
            .I(N__40353));
    Span4Mux_v I__8578 (
            .O(N__40353),
            .I(N__40350));
    Odrv4 I__8577 (
            .O(N__40350),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__8576 (
            .O(N__40347),
            .I(N__40344));
    LocalMux I__8575 (
            .O(N__40344),
            .I(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ));
    InMux I__8574 (
            .O(N__40341),
            .I(N__40338));
    LocalMux I__8573 (
            .O(N__40338),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__8572 (
            .O(N__40335),
            .I(N__40332));
    LocalMux I__8571 (
            .O(N__40332),
            .I(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ));
    CascadeMux I__8570 (
            .O(N__40329),
            .I(N__40326));
    InMux I__8569 (
            .O(N__40326),
            .I(N__40323));
    LocalMux I__8568 (
            .O(N__40323),
            .I(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ));
    InMux I__8567 (
            .O(N__40320),
            .I(N__40315));
    InMux I__8566 (
            .O(N__40319),
            .I(N__40311));
    InMux I__8565 (
            .O(N__40318),
            .I(N__40308));
    LocalMux I__8564 (
            .O(N__40315),
            .I(N__40305));
    InMux I__8563 (
            .O(N__40314),
            .I(N__40302));
    LocalMux I__8562 (
            .O(N__40311),
            .I(N__40297));
    LocalMux I__8561 (
            .O(N__40308),
            .I(N__40297));
    Span4Mux_h I__8560 (
            .O(N__40305),
            .I(N__40294));
    LocalMux I__8559 (
            .O(N__40302),
            .I(N__40291));
    Span4Mux_h I__8558 (
            .O(N__40297),
            .I(N__40288));
    Span4Mux_h I__8557 (
            .O(N__40294),
            .I(N__40285));
    Odrv12 I__8556 (
            .O(N__40291),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__8555 (
            .O(N__40288),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__8554 (
            .O(N__40285),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__8553 (
            .O(N__40278),
            .I(N__40275));
    InMux I__8552 (
            .O(N__40275),
            .I(N__40272));
    LocalMux I__8551 (
            .O(N__40272),
            .I(N__40269));
    Span4Mux_h I__8550 (
            .O(N__40269),
            .I(N__40266));
    Span4Mux_h I__8549 (
            .O(N__40266),
            .I(N__40263));
    Odrv4 I__8548 (
            .O(N__40263),
            .I(\current_shift_inst.PI_CTRL.integrator_i_29 ));
    InMux I__8547 (
            .O(N__40260),
            .I(N__40257));
    LocalMux I__8546 (
            .O(N__40257),
            .I(N__40253));
    InMux I__8545 (
            .O(N__40256),
            .I(N__40250));
    Span4Mux_v I__8544 (
            .O(N__40253),
            .I(N__40245));
    LocalMux I__8543 (
            .O(N__40250),
            .I(N__40245));
    Span4Mux_v I__8542 (
            .O(N__40245),
            .I(N__40240));
    InMux I__8541 (
            .O(N__40244),
            .I(N__40235));
    InMux I__8540 (
            .O(N__40243),
            .I(N__40235));
    Odrv4 I__8539 (
            .O(N__40240),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__8538 (
            .O(N__40235),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__8537 (
            .O(N__40230),
            .I(N__40227));
    LocalMux I__8536 (
            .O(N__40227),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__8535 (
            .O(N__40224),
            .I(N__40219));
    InMux I__8534 (
            .O(N__40223),
            .I(N__40216));
    InMux I__8533 (
            .O(N__40222),
            .I(N__40213));
    LocalMux I__8532 (
            .O(N__40219),
            .I(N__40208));
    LocalMux I__8531 (
            .O(N__40216),
            .I(N__40208));
    LocalMux I__8530 (
            .O(N__40213),
            .I(N__40205));
    Span4Mux_v I__8529 (
            .O(N__40208),
            .I(N__40201));
    Span4Mux_h I__8528 (
            .O(N__40205),
            .I(N__40198));
    InMux I__8527 (
            .O(N__40204),
            .I(N__40195));
    Odrv4 I__8526 (
            .O(N__40201),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__8525 (
            .O(N__40198),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__8524 (
            .O(N__40195),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    CascadeMux I__8523 (
            .O(N__40188),
            .I(N__40185));
    InMux I__8522 (
            .O(N__40185),
            .I(N__40182));
    LocalMux I__8521 (
            .O(N__40182),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    CascadeMux I__8520 (
            .O(N__40179),
            .I(N__40176));
    InMux I__8519 (
            .O(N__40176),
            .I(N__40173));
    LocalMux I__8518 (
            .O(N__40173),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    CascadeMux I__8517 (
            .O(N__40170),
            .I(N__40167));
    InMux I__8516 (
            .O(N__40167),
            .I(N__40164));
    LocalMux I__8515 (
            .O(N__40164),
            .I(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ));
    InMux I__8514 (
            .O(N__40161),
            .I(N__40158));
    LocalMux I__8513 (
            .O(N__40158),
            .I(N__40155));
    Span4Mux_h I__8512 (
            .O(N__40155),
            .I(N__40152));
    Odrv4 I__8511 (
            .O(N__40152),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__8510 (
            .O(N__40149),
            .I(N__40146));
    LocalMux I__8509 (
            .O(N__40146),
            .I(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ));
    CascadeMux I__8508 (
            .O(N__40143),
            .I(N__40140));
    InMux I__8507 (
            .O(N__40140),
            .I(N__40137));
    LocalMux I__8506 (
            .O(N__40137),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    CascadeMux I__8505 (
            .O(N__40134),
            .I(N__40131));
    InMux I__8504 (
            .O(N__40131),
            .I(N__40127));
    CascadeMux I__8503 (
            .O(N__40130),
            .I(N__40124));
    LocalMux I__8502 (
            .O(N__40127),
            .I(N__40120));
    InMux I__8501 (
            .O(N__40124),
            .I(N__40117));
    InMux I__8500 (
            .O(N__40123),
            .I(N__40114));
    Span4Mux_v I__8499 (
            .O(N__40120),
            .I(N__40110));
    LocalMux I__8498 (
            .O(N__40117),
            .I(N__40107));
    LocalMux I__8497 (
            .O(N__40114),
            .I(N__40104));
    InMux I__8496 (
            .O(N__40113),
            .I(N__40101));
    Span4Mux_v I__8495 (
            .O(N__40110),
            .I(N__40092));
    Span4Mux_v I__8494 (
            .O(N__40107),
            .I(N__40092));
    Span4Mux_h I__8493 (
            .O(N__40104),
            .I(N__40092));
    LocalMux I__8492 (
            .O(N__40101),
            .I(N__40092));
    Odrv4 I__8491 (
            .O(N__40092),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__8490 (
            .O(N__40089),
            .I(N__40086));
    LocalMux I__8489 (
            .O(N__40086),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    CascadeMux I__8488 (
            .O(N__40083),
            .I(N__40080));
    InMux I__8487 (
            .O(N__40080),
            .I(N__40077));
    LocalMux I__8486 (
            .O(N__40077),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    CascadeMux I__8485 (
            .O(N__40074),
            .I(N__40069));
    CascadeMux I__8484 (
            .O(N__40073),
            .I(N__40066));
    InMux I__8483 (
            .O(N__40072),
            .I(N__40063));
    InMux I__8482 (
            .O(N__40069),
            .I(N__40059));
    InMux I__8481 (
            .O(N__40066),
            .I(N__40056));
    LocalMux I__8480 (
            .O(N__40063),
            .I(N__40053));
    CascadeMux I__8479 (
            .O(N__40062),
            .I(N__40050));
    LocalMux I__8478 (
            .O(N__40059),
            .I(N__40046));
    LocalMux I__8477 (
            .O(N__40056),
            .I(N__40043));
    Span4Mux_h I__8476 (
            .O(N__40053),
            .I(N__40040));
    InMux I__8475 (
            .O(N__40050),
            .I(N__40035));
    InMux I__8474 (
            .O(N__40049),
            .I(N__40035));
    Span4Mux_h I__8473 (
            .O(N__40046),
            .I(N__40030));
    Span4Mux_v I__8472 (
            .O(N__40043),
            .I(N__40030));
    Span4Mux_h I__8471 (
            .O(N__40040),
            .I(N__40027));
    LocalMux I__8470 (
            .O(N__40035),
            .I(N__40024));
    Odrv4 I__8469 (
            .O(N__40030),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__8468 (
            .O(N__40027),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__8467 (
            .O(N__40024),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__8466 (
            .O(N__40017),
            .I(N__40014));
    LocalMux I__8465 (
            .O(N__40014),
            .I(N__40011));
    Span4Mux_v I__8464 (
            .O(N__40011),
            .I(N__40008));
    Span4Mux_h I__8463 (
            .O(N__40008),
            .I(N__40005));
    Odrv4 I__8462 (
            .O(N__40005),
            .I(\current_shift_inst.PI_CTRL.integrator_i_26 ));
    CascadeMux I__8461 (
            .O(N__40002),
            .I(N__39999));
    InMux I__8460 (
            .O(N__39999),
            .I(N__39996));
    LocalMux I__8459 (
            .O(N__39996),
            .I(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ));
    InMux I__8458 (
            .O(N__39993),
            .I(N__39990));
    LocalMux I__8457 (
            .O(N__39990),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__8456 (
            .O(N__39987),
            .I(N__39984));
    LocalMux I__8455 (
            .O(N__39984),
            .I(N__39981));
    Span4Mux_v I__8454 (
            .O(N__39981),
            .I(N__39977));
    InMux I__8453 (
            .O(N__39980),
            .I(N__39974));
    Sp12to4 I__8452 (
            .O(N__39977),
            .I(N__39968));
    LocalMux I__8451 (
            .O(N__39974),
            .I(N__39968));
    InMux I__8450 (
            .O(N__39973),
            .I(N__39965));
    Odrv12 I__8449 (
            .O(N__39968),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    LocalMux I__8448 (
            .O(N__39965),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CascadeMux I__8447 (
            .O(N__39960),
            .I(N__39957));
    InMux I__8446 (
            .O(N__39957),
            .I(N__39954));
    LocalMux I__8445 (
            .O(N__39954),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    CascadeMux I__8444 (
            .O(N__39951),
            .I(N__39948));
    InMux I__8443 (
            .O(N__39948),
            .I(N__39942));
    InMux I__8442 (
            .O(N__39947),
            .I(N__39942));
    LocalMux I__8441 (
            .O(N__39942),
            .I(N__39937));
    InMux I__8440 (
            .O(N__39941),
            .I(N__39932));
    InMux I__8439 (
            .O(N__39940),
            .I(N__39932));
    Span4Mux_v I__8438 (
            .O(N__39937),
            .I(N__39927));
    LocalMux I__8437 (
            .O(N__39932),
            .I(N__39927));
    Odrv4 I__8436 (
            .O(N__39927),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    CascadeMux I__8435 (
            .O(N__39924),
            .I(N__39921));
    InMux I__8434 (
            .O(N__39921),
            .I(N__39918));
    LocalMux I__8433 (
            .O(N__39918),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    InMux I__8432 (
            .O(N__39915),
            .I(N__39912));
    LocalMux I__8431 (
            .O(N__39912),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__8430 (
            .O(N__39909),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    CascadeMux I__8429 (
            .O(N__39906),
            .I(N__39903));
    InMux I__8428 (
            .O(N__39903),
            .I(N__39900));
    LocalMux I__8427 (
            .O(N__39900),
            .I(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ));
    CascadeMux I__8426 (
            .O(N__39897),
            .I(N__39894));
    InMux I__8425 (
            .O(N__39894),
            .I(N__39891));
    LocalMux I__8424 (
            .O(N__39891),
            .I(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ));
    InMux I__8423 (
            .O(N__39888),
            .I(N__39885));
    LocalMux I__8422 (
            .O(N__39885),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__8421 (
            .O(N__39882),
            .I(N__39879));
    InMux I__8420 (
            .O(N__39879),
            .I(N__39876));
    LocalMux I__8419 (
            .O(N__39876),
            .I(N__39873));
    Span4Mux_h I__8418 (
            .O(N__39873),
            .I(N__39870));
    Span4Mux_v I__8417 (
            .O(N__39870),
            .I(N__39867));
    Odrv4 I__8416 (
            .O(N__39867),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    CascadeMux I__8415 (
            .O(N__39864),
            .I(N__39860));
    InMux I__8414 (
            .O(N__39863),
            .I(N__39852));
    InMux I__8413 (
            .O(N__39860),
            .I(N__39852));
    InMux I__8412 (
            .O(N__39859),
            .I(N__39852));
    LocalMux I__8411 (
            .O(N__39852),
            .I(N__39848));
    InMux I__8410 (
            .O(N__39851),
            .I(N__39845));
    Odrv4 I__8409 (
            .O(N__39848),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__8408 (
            .O(N__39845),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    CascadeMux I__8407 (
            .O(N__39840),
            .I(N__39837));
    InMux I__8406 (
            .O(N__39837),
            .I(N__39834));
    LocalMux I__8405 (
            .O(N__39834),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__8404 (
            .O(N__39831),
            .I(N__39828));
    LocalMux I__8403 (
            .O(N__39828),
            .I(N__39825));
    Span4Mux_v I__8402 (
            .O(N__39825),
            .I(N__39822));
    Odrv4 I__8401 (
            .O(N__39822),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__8400 (
            .O(N__39819),
            .I(N__39816));
    LocalMux I__8399 (
            .O(N__39816),
            .I(N__39813));
    Span4Mux_v I__8398 (
            .O(N__39813),
            .I(N__39810));
    Odrv4 I__8397 (
            .O(N__39810),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    CascadeMux I__8396 (
            .O(N__39807),
            .I(N__39803));
    InMux I__8395 (
            .O(N__39806),
            .I(N__39795));
    InMux I__8394 (
            .O(N__39803),
            .I(N__39795));
    InMux I__8393 (
            .O(N__39802),
            .I(N__39795));
    LocalMux I__8392 (
            .O(N__39795),
            .I(N__39792));
    Span4Mux_h I__8391 (
            .O(N__39792),
            .I(N__39788));
    InMux I__8390 (
            .O(N__39791),
            .I(N__39785));
    Odrv4 I__8389 (
            .O(N__39788),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__8388 (
            .O(N__39785),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__8387 (
            .O(N__39780),
            .I(N__39777));
    LocalMux I__8386 (
            .O(N__39777),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__8385 (
            .O(N__39774),
            .I(N__39771));
    InMux I__8384 (
            .O(N__39771),
            .I(N__39768));
    LocalMux I__8383 (
            .O(N__39768),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    CascadeMux I__8382 (
            .O(N__39765),
            .I(N__39762));
    InMux I__8381 (
            .O(N__39762),
            .I(N__39759));
    LocalMux I__8380 (
            .O(N__39759),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    CascadeMux I__8379 (
            .O(N__39756),
            .I(N__39753));
    InMux I__8378 (
            .O(N__39753),
            .I(N__39750));
    LocalMux I__8377 (
            .O(N__39750),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    CascadeMux I__8376 (
            .O(N__39747),
            .I(N__39744));
    InMux I__8375 (
            .O(N__39744),
            .I(N__39741));
    LocalMux I__8374 (
            .O(N__39741),
            .I(N__39738));
    Span4Mux_v I__8373 (
            .O(N__39738),
            .I(N__39735));
    Odrv4 I__8372 (
            .O(N__39735),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    CascadeMux I__8371 (
            .O(N__39732),
            .I(N__39729));
    InMux I__8370 (
            .O(N__39729),
            .I(N__39726));
    LocalMux I__8369 (
            .O(N__39726),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    CascadeMux I__8368 (
            .O(N__39723),
            .I(N__39720));
    InMux I__8367 (
            .O(N__39720),
            .I(N__39717));
    LocalMux I__8366 (
            .O(N__39717),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    InMux I__8365 (
            .O(N__39714),
            .I(N__39711));
    LocalMux I__8364 (
            .O(N__39711),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    InMux I__8363 (
            .O(N__39708),
            .I(N__39705));
    LocalMux I__8362 (
            .O(N__39705),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__8361 (
            .O(N__39702),
            .I(N__39699));
    LocalMux I__8360 (
            .O(N__39699),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__8359 (
            .O(N__39696),
            .I(N__39693));
    LocalMux I__8358 (
            .O(N__39693),
            .I(N__39690));
    Span12Mux_h I__8357 (
            .O(N__39690),
            .I(N__39687));
    Odrv12 I__8356 (
            .O(N__39687),
            .I(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ));
    CascadeMux I__8355 (
            .O(N__39684),
            .I(N__39678));
    InMux I__8354 (
            .O(N__39683),
            .I(N__39673));
    InMux I__8353 (
            .O(N__39682),
            .I(N__39673));
    InMux I__8352 (
            .O(N__39681),
            .I(N__39668));
    InMux I__8351 (
            .O(N__39678),
            .I(N__39668));
    LocalMux I__8350 (
            .O(N__39673),
            .I(N__39665));
    LocalMux I__8349 (
            .O(N__39668),
            .I(N__39662));
    Span4Mux_v I__8348 (
            .O(N__39665),
            .I(N__39659));
    Odrv12 I__8347 (
            .O(N__39662),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv4 I__8346 (
            .O(N__39659),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    CascadeMux I__8345 (
            .O(N__39654),
            .I(N__39651));
    InMux I__8344 (
            .O(N__39651),
            .I(N__39648));
    LocalMux I__8343 (
            .O(N__39648),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    CascadeMux I__8342 (
            .O(N__39645),
            .I(N__39642));
    InMux I__8341 (
            .O(N__39642),
            .I(N__39639));
    LocalMux I__8340 (
            .O(N__39639),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__8339 (
            .O(N__39636),
            .I(N__39633));
    LocalMux I__8338 (
            .O(N__39633),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    InMux I__8337 (
            .O(N__39630),
            .I(N__39627));
    LocalMux I__8336 (
            .O(N__39627),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__8335 (
            .O(N__39624),
            .I(N__39621));
    InMux I__8334 (
            .O(N__39621),
            .I(N__39618));
    LocalMux I__8333 (
            .O(N__39618),
            .I(N__39615));
    Odrv4 I__8332 (
            .O(N__39615),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__8331 (
            .O(N__39612),
            .I(N__39608));
    InMux I__8330 (
            .O(N__39611),
            .I(N__39605));
    LocalMux I__8329 (
            .O(N__39608),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__8328 (
            .O(N__39605),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__8327 (
            .O(N__39600),
            .I(N__39596));
    InMux I__8326 (
            .O(N__39599),
            .I(N__39593));
    LocalMux I__8325 (
            .O(N__39596),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__8324 (
            .O(N__39593),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__8323 (
            .O(N__39588),
            .I(N__39585));
    LocalMux I__8322 (
            .O(N__39585),
            .I(N__39582));
    Odrv4 I__8321 (
            .O(N__39582),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df26 ));
    InMux I__8320 (
            .O(N__39579),
            .I(N__39574));
    InMux I__8319 (
            .O(N__39578),
            .I(N__39571));
    InMux I__8318 (
            .O(N__39577),
            .I(N__39568));
    LocalMux I__8317 (
            .O(N__39574),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__8316 (
            .O(N__39571),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__8315 (
            .O(N__39568),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__8314 (
            .O(N__39561),
            .I(N__39556));
    InMux I__8313 (
            .O(N__39560),
            .I(N__39553));
    InMux I__8312 (
            .O(N__39559),
            .I(N__39550));
    LocalMux I__8311 (
            .O(N__39556),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__8310 (
            .O(N__39553),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__8309 (
            .O(N__39550),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    CascadeMux I__8308 (
            .O(N__39543),
            .I(N__39540));
    InMux I__8307 (
            .O(N__39540),
            .I(N__39537));
    LocalMux I__8306 (
            .O(N__39537),
            .I(N__39534));
    Odrv4 I__8305 (
            .O(N__39534),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__8304 (
            .O(N__39531),
            .I(N__39528));
    LocalMux I__8303 (
            .O(N__39528),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    InMux I__8302 (
            .O(N__39525),
            .I(N__39520));
    InMux I__8301 (
            .O(N__39524),
            .I(N__39515));
    InMux I__8300 (
            .O(N__39523),
            .I(N__39515));
    LocalMux I__8299 (
            .O(N__39520),
            .I(N__39511));
    LocalMux I__8298 (
            .O(N__39515),
            .I(N__39508));
    InMux I__8297 (
            .O(N__39514),
            .I(N__39505));
    Span4Mux_v I__8296 (
            .O(N__39511),
            .I(N__39498));
    Span4Mux_h I__8295 (
            .O(N__39508),
            .I(N__39498));
    LocalMux I__8294 (
            .O(N__39505),
            .I(N__39498));
    Odrv4 I__8293 (
            .O(N__39498),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__8292 (
            .O(N__39495),
            .I(N__39492));
    LocalMux I__8291 (
            .O(N__39492),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__8290 (
            .O(N__39489),
            .I(N__39486));
    InMux I__8289 (
            .O(N__39486),
            .I(N__39483));
    LocalMux I__8288 (
            .O(N__39483),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    CascadeMux I__8287 (
            .O(N__39480),
            .I(N__39477));
    InMux I__8286 (
            .O(N__39477),
            .I(N__39474));
    LocalMux I__8285 (
            .O(N__39474),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__8284 (
            .O(N__39471),
            .I(N__39468));
    LocalMux I__8283 (
            .O(N__39468),
            .I(N__39465));
    Odrv4 I__8282 (
            .O(N__39465),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ));
    InMux I__8281 (
            .O(N__39462),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ));
    InMux I__8280 (
            .O(N__39459),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    InMux I__8279 (
            .O(N__39456),
            .I(N__39452));
    InMux I__8278 (
            .O(N__39455),
            .I(N__39449));
    LocalMux I__8277 (
            .O(N__39452),
            .I(N__39446));
    LocalMux I__8276 (
            .O(N__39449),
            .I(N__39443));
    Span4Mux_h I__8275 (
            .O(N__39446),
            .I(N__39440));
    Odrv4 I__8274 (
            .O(N__39443),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__8273 (
            .O(N__39440),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__8272 (
            .O(N__39435),
            .I(N__39432));
    LocalMux I__8271 (
            .O(N__39432),
            .I(N__39429));
    Odrv4 I__8270 (
            .O(N__39429),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    InMux I__8269 (
            .O(N__39426),
            .I(N__39419));
    InMux I__8268 (
            .O(N__39425),
            .I(N__39419));
    InMux I__8267 (
            .O(N__39424),
            .I(N__39416));
    LocalMux I__8266 (
            .O(N__39419),
            .I(N__39413));
    LocalMux I__8265 (
            .O(N__39416),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__8264 (
            .O(N__39413),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__8263 (
            .O(N__39408),
            .I(N__39403));
    InMux I__8262 (
            .O(N__39407),
            .I(N__39398));
    InMux I__8261 (
            .O(N__39406),
            .I(N__39398));
    LocalMux I__8260 (
            .O(N__39403),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__8259 (
            .O(N__39398),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__8258 (
            .O(N__39393),
            .I(N__39390));
    InMux I__8257 (
            .O(N__39390),
            .I(N__39387));
    LocalMux I__8256 (
            .O(N__39387),
            .I(N__39384));
    Span4Mux_h I__8255 (
            .O(N__39384),
            .I(N__39381));
    Odrv4 I__8254 (
            .O(N__39381),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    CascadeMux I__8253 (
            .O(N__39378),
            .I(N__39375));
    InMux I__8252 (
            .O(N__39375),
            .I(N__39369));
    InMux I__8251 (
            .O(N__39374),
            .I(N__39369));
    LocalMux I__8250 (
            .O(N__39369),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__8249 (
            .O(N__39366),
            .I(N__39363));
    LocalMux I__8248 (
            .O(N__39363),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    InMux I__8247 (
            .O(N__39360),
            .I(N__39355));
    InMux I__8246 (
            .O(N__39359),
            .I(N__39351));
    InMux I__8245 (
            .O(N__39358),
            .I(N__39348));
    LocalMux I__8244 (
            .O(N__39355),
            .I(N__39345));
    InMux I__8243 (
            .O(N__39354),
            .I(N__39342));
    LocalMux I__8242 (
            .O(N__39351),
            .I(N__39339));
    LocalMux I__8241 (
            .O(N__39348),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__8240 (
            .O(N__39345),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__8239 (
            .O(N__39342),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv12 I__8238 (
            .O(N__39339),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    CascadeMux I__8237 (
            .O(N__39330),
            .I(N__39327));
    InMux I__8236 (
            .O(N__39327),
            .I(N__39324));
    LocalMux I__8235 (
            .O(N__39324),
            .I(N__39319));
    InMux I__8234 (
            .O(N__39323),
            .I(N__39316));
    InMux I__8233 (
            .O(N__39322),
            .I(N__39313));
    Span4Mux_h I__8232 (
            .O(N__39319),
            .I(N__39310));
    LocalMux I__8231 (
            .O(N__39316),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__8230 (
            .O(N__39313),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__8229 (
            .O(N__39310),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    CascadeMux I__8228 (
            .O(N__39303),
            .I(N__39300));
    InMux I__8227 (
            .O(N__39300),
            .I(N__39297));
    LocalMux I__8226 (
            .O(N__39297),
            .I(N__39294));
    Odrv4 I__8225 (
            .O(N__39294),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ));
    InMux I__8224 (
            .O(N__39291),
            .I(N__39287));
    InMux I__8223 (
            .O(N__39290),
            .I(N__39284));
    LocalMux I__8222 (
            .O(N__39287),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__8221 (
            .O(N__39284),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__8220 (
            .O(N__39279),
            .I(N__39275));
    InMux I__8219 (
            .O(N__39278),
            .I(N__39272));
    LocalMux I__8218 (
            .O(N__39275),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__8217 (
            .O(N__39272),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__8216 (
            .O(N__39267),
            .I(N__39264));
    LocalMux I__8215 (
            .O(N__39264),
            .I(N__39261));
    Odrv12 I__8214 (
            .O(N__39261),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df28 ));
    InMux I__8213 (
            .O(N__39258),
            .I(N__39255));
    LocalMux I__8212 (
            .O(N__39255),
            .I(N__39252));
    Odrv4 I__8211 (
            .O(N__39252),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__8210 (
            .O(N__39249),
            .I(N__39245));
    InMux I__8209 (
            .O(N__39248),
            .I(N__39242));
    LocalMux I__8208 (
            .O(N__39245),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__8207 (
            .O(N__39242),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__8206 (
            .O(N__39237),
            .I(N__39234));
    InMux I__8205 (
            .O(N__39234),
            .I(N__39231));
    LocalMux I__8204 (
            .O(N__39231),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__8203 (
            .O(N__39228),
            .I(N__39225));
    InMux I__8202 (
            .O(N__39225),
            .I(N__39222));
    LocalMux I__8201 (
            .O(N__39222),
            .I(N__39219));
    Odrv12 I__8200 (
            .O(N__39219),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__8199 (
            .O(N__39216),
            .I(N__39212));
    InMux I__8198 (
            .O(N__39215),
            .I(N__39209));
    LocalMux I__8197 (
            .O(N__39212),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__8196 (
            .O(N__39209),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__8195 (
            .O(N__39204),
            .I(N__39201));
    LocalMux I__8194 (
            .O(N__39201),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__8193 (
            .O(N__39198),
            .I(N__39195));
    LocalMux I__8192 (
            .O(N__39195),
            .I(N__39192));
    Odrv4 I__8191 (
            .O(N__39192),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df20 ));
    InMux I__8190 (
            .O(N__39189),
            .I(N__39186));
    LocalMux I__8189 (
            .O(N__39186),
            .I(N__39183));
    Span4Mux_v I__8188 (
            .O(N__39183),
            .I(N__39180));
    Odrv4 I__8187 (
            .O(N__39180),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df22 ));
    InMux I__8186 (
            .O(N__39177),
            .I(N__39174));
    LocalMux I__8185 (
            .O(N__39174),
            .I(N__39171));
    Odrv4 I__8184 (
            .O(N__39171),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df24 ));
    InMux I__8183 (
            .O(N__39168),
            .I(N__39164));
    InMux I__8182 (
            .O(N__39167),
            .I(N__39161));
    LocalMux I__8181 (
            .O(N__39164),
            .I(N__39158));
    LocalMux I__8180 (
            .O(N__39161),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__8179 (
            .O(N__39158),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__8178 (
            .O(N__39153),
            .I(N__39150));
    InMux I__8177 (
            .O(N__39150),
            .I(N__39147));
    LocalMux I__8176 (
            .O(N__39147),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__8175 (
            .O(N__39144),
            .I(N__39141));
    InMux I__8174 (
            .O(N__39141),
            .I(N__39138));
    LocalMux I__8173 (
            .O(N__39138),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    InMux I__8172 (
            .O(N__39135),
            .I(N__39131));
    InMux I__8171 (
            .O(N__39134),
            .I(N__39128));
    LocalMux I__8170 (
            .O(N__39131),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__8169 (
            .O(N__39128),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__8168 (
            .O(N__39123),
            .I(N__39120));
    LocalMux I__8167 (
            .O(N__39120),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__8166 (
            .O(N__39117),
            .I(N__39113));
    InMux I__8165 (
            .O(N__39116),
            .I(N__39110));
    LocalMux I__8164 (
            .O(N__39113),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__8163 (
            .O(N__39110),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__8162 (
            .O(N__39105),
            .I(N__39102));
    InMux I__8161 (
            .O(N__39102),
            .I(N__39099));
    LocalMux I__8160 (
            .O(N__39099),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    InMux I__8159 (
            .O(N__39096),
            .I(N__39093));
    LocalMux I__8158 (
            .O(N__39093),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__8157 (
            .O(N__39090),
            .I(N__39086));
    InMux I__8156 (
            .O(N__39089),
            .I(N__39083));
    LocalMux I__8155 (
            .O(N__39086),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__8154 (
            .O(N__39083),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    CascadeMux I__8153 (
            .O(N__39078),
            .I(N__39075));
    InMux I__8152 (
            .O(N__39075),
            .I(N__39072));
    LocalMux I__8151 (
            .O(N__39072),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__8150 (
            .O(N__39069),
            .I(N__39065));
    InMux I__8149 (
            .O(N__39068),
            .I(N__39062));
    LocalMux I__8148 (
            .O(N__39065),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__8147 (
            .O(N__39062),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__8146 (
            .O(N__39057),
            .I(N__39054));
    LocalMux I__8145 (
            .O(N__39054),
            .I(N__39051));
    Span4Mux_h I__8144 (
            .O(N__39051),
            .I(N__39048));
    Odrv4 I__8143 (
            .O(N__39048),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__8142 (
            .O(N__39045),
            .I(N__39042));
    InMux I__8141 (
            .O(N__39042),
            .I(N__39039));
    LocalMux I__8140 (
            .O(N__39039),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__8139 (
            .O(N__39036),
            .I(N__39033));
    LocalMux I__8138 (
            .O(N__39033),
            .I(N__39030));
    Span4Mux_v I__8137 (
            .O(N__39030),
            .I(N__39027));
    Span4Mux_v I__8136 (
            .O(N__39027),
            .I(N__39024));
    Odrv4 I__8135 (
            .O(N__39024),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__8134 (
            .O(N__39021),
            .I(N__39017));
    InMux I__8133 (
            .O(N__39020),
            .I(N__39014));
    LocalMux I__8132 (
            .O(N__39017),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__8131 (
            .O(N__39014),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    CascadeMux I__8130 (
            .O(N__39009),
            .I(N__39006));
    InMux I__8129 (
            .O(N__39006),
            .I(N__39003));
    LocalMux I__8128 (
            .O(N__39003),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__8127 (
            .O(N__39000),
            .I(N__38996));
    InMux I__8126 (
            .O(N__38999),
            .I(N__38993));
    LocalMux I__8125 (
            .O(N__38996),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__8124 (
            .O(N__38993),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    CascadeMux I__8123 (
            .O(N__38988),
            .I(N__38985));
    InMux I__8122 (
            .O(N__38985),
            .I(N__38982));
    LocalMux I__8121 (
            .O(N__38982),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__8120 (
            .O(N__38979),
            .I(N__38975));
    InMux I__8119 (
            .O(N__38978),
            .I(N__38972));
    LocalMux I__8118 (
            .O(N__38975),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__8117 (
            .O(N__38972),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__8116 (
            .O(N__38967),
            .I(N__38964));
    InMux I__8115 (
            .O(N__38964),
            .I(N__38961));
    LocalMux I__8114 (
            .O(N__38961),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__8113 (
            .O(N__38958),
            .I(N__38954));
    CascadeMux I__8112 (
            .O(N__38957),
            .I(N__38951));
    InMux I__8111 (
            .O(N__38954),
            .I(N__38948));
    InMux I__8110 (
            .O(N__38951),
            .I(N__38944));
    LocalMux I__8109 (
            .O(N__38948),
            .I(N__38941));
    InMux I__8108 (
            .O(N__38947),
            .I(N__38938));
    LocalMux I__8107 (
            .O(N__38944),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__8106 (
            .O(N__38941),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__8105 (
            .O(N__38938),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__8104 (
            .O(N__38931),
            .I(N__38928));
    InMux I__8103 (
            .O(N__38928),
            .I(N__38925));
    LocalMux I__8102 (
            .O(N__38925),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__8101 (
            .O(N__38922),
            .I(N__38918));
    InMux I__8100 (
            .O(N__38921),
            .I(N__38915));
    LocalMux I__8099 (
            .O(N__38918),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__8098 (
            .O(N__38915),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    CascadeMux I__8097 (
            .O(N__38910),
            .I(N__38907));
    InMux I__8096 (
            .O(N__38907),
            .I(N__38904));
    LocalMux I__8095 (
            .O(N__38904),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__8094 (
            .O(N__38901),
            .I(N__38897));
    InMux I__8093 (
            .O(N__38900),
            .I(N__38894));
    LocalMux I__8092 (
            .O(N__38897),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__8091 (
            .O(N__38894),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__8090 (
            .O(N__38889),
            .I(N__38886));
    InMux I__8089 (
            .O(N__38886),
            .I(N__38883));
    LocalMux I__8088 (
            .O(N__38883),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__8087 (
            .O(N__38880),
            .I(N__38876));
    InMux I__8086 (
            .O(N__38879),
            .I(N__38873));
    LocalMux I__8085 (
            .O(N__38876),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__8084 (
            .O(N__38873),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__8083 (
            .O(N__38868),
            .I(N__38865));
    InMux I__8082 (
            .O(N__38865),
            .I(N__38862));
    LocalMux I__8081 (
            .O(N__38862),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__8080 (
            .O(N__38859),
            .I(N__38855));
    InMux I__8079 (
            .O(N__38858),
            .I(N__38852));
    LocalMux I__8078 (
            .O(N__38855),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__8077 (
            .O(N__38852),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__8076 (
            .O(N__38847),
            .I(N__38844));
    LocalMux I__8075 (
            .O(N__38844),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__8074 (
            .O(N__38841),
            .I(N__38838));
    InMux I__8073 (
            .O(N__38838),
            .I(N__38835));
    LocalMux I__8072 (
            .O(N__38835),
            .I(N__38832));
    Odrv4 I__8071 (
            .O(N__38832),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__8070 (
            .O(N__38829),
            .I(N__38826));
    LocalMux I__8069 (
            .O(N__38826),
            .I(N__38823));
    Span4Mux_h I__8068 (
            .O(N__38823),
            .I(N__38820));
    Span4Mux_h I__8067 (
            .O(N__38820),
            .I(N__38817));
    Odrv4 I__8066 (
            .O(N__38817),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    InMux I__8065 (
            .O(N__38814),
            .I(N__38807));
    InMux I__8064 (
            .O(N__38813),
            .I(N__38807));
    InMux I__8063 (
            .O(N__38812),
            .I(N__38804));
    LocalMux I__8062 (
            .O(N__38807),
            .I(N__38801));
    LocalMux I__8061 (
            .O(N__38804),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__8060 (
            .O(N__38801),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__8059 (
            .O(N__38796),
            .I(N__38793));
    InMux I__8058 (
            .O(N__38793),
            .I(N__38787));
    InMux I__8057 (
            .O(N__38792),
            .I(N__38787));
    LocalMux I__8056 (
            .O(N__38787),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    InMux I__8055 (
            .O(N__38784),
            .I(N__38779));
    InMux I__8054 (
            .O(N__38783),
            .I(N__38774));
    InMux I__8053 (
            .O(N__38782),
            .I(N__38774));
    LocalMux I__8052 (
            .O(N__38779),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__8051 (
            .O(N__38774),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__8050 (
            .O(N__38769),
            .I(N__38766));
    InMux I__8049 (
            .O(N__38766),
            .I(N__38763));
    LocalMux I__8048 (
            .O(N__38763),
            .I(N__38760));
    Odrv12 I__8047 (
            .O(N__38760),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    CascadeMux I__8046 (
            .O(N__38757),
            .I(elapsed_time_ns_1_RNIQENQL1_0_9_cascade_));
    InMux I__8045 (
            .O(N__38754),
            .I(N__38751));
    LocalMux I__8044 (
            .O(N__38751),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ));
    CascadeMux I__8043 (
            .O(N__38748),
            .I(\phase_controller_inst1.stoper_tr.N_242_cascade_ ));
    InMux I__8042 (
            .O(N__38745),
            .I(N__38742));
    LocalMux I__8041 (
            .O(N__38742),
            .I(N__38739));
    Span4Mux_h I__8040 (
            .O(N__38739),
            .I(N__38736));
    Odrv4 I__8039 (
            .O(N__38736),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    InMux I__8038 (
            .O(N__38733),
            .I(N__38730));
    LocalMux I__8037 (
            .O(N__38730),
            .I(N__38727));
    Span4Mux_v I__8036 (
            .O(N__38727),
            .I(N__38724));
    Span4Mux_h I__8035 (
            .O(N__38724),
            .I(N__38721));
    Sp12to4 I__8034 (
            .O(N__38721),
            .I(N__38718));
    Odrv12 I__8033 (
            .O(N__38718),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    InMux I__8032 (
            .O(N__38715),
            .I(N__38712));
    LocalMux I__8031 (
            .O(N__38712),
            .I(N__38709));
    Span4Mux_h I__8030 (
            .O(N__38709),
            .I(N__38706));
    Odrv4 I__8029 (
            .O(N__38706),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9 ));
    CascadeMux I__8028 (
            .O(N__38703),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ));
    InMux I__8027 (
            .O(N__38700),
            .I(N__38697));
    LocalMux I__8026 (
            .O(N__38697),
            .I(N__38694));
    Span4Mux_h I__8025 (
            .O(N__38694),
            .I(N__38691));
    Odrv4 I__8024 (
            .O(N__38691),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    InMux I__8023 (
            .O(N__38688),
            .I(N__38685));
    LocalMux I__8022 (
            .O(N__38685),
            .I(N__38682));
    Span4Mux_h I__8021 (
            .O(N__38682),
            .I(N__38679));
    Odrv4 I__8020 (
            .O(N__38679),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    CascadeMux I__8019 (
            .O(N__38676),
            .I(N__38673));
    InMux I__8018 (
            .O(N__38673),
            .I(N__38669));
    InMux I__8017 (
            .O(N__38672),
            .I(N__38666));
    LocalMux I__8016 (
            .O(N__38669),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    LocalMux I__8015 (
            .O(N__38666),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    CascadeMux I__8014 (
            .O(N__38661),
            .I(N__38656));
    InMux I__8013 (
            .O(N__38660),
            .I(N__38653));
    InMux I__8012 (
            .O(N__38659),
            .I(N__38648));
    InMux I__8011 (
            .O(N__38656),
            .I(N__38648));
    LocalMux I__8010 (
            .O(N__38653),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__8009 (
            .O(N__38648),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__8008 (
            .O(N__38643),
            .I(N__38638));
    InMux I__8007 (
            .O(N__38642),
            .I(N__38635));
    InMux I__8006 (
            .O(N__38641),
            .I(N__38632));
    LocalMux I__8005 (
            .O(N__38638),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__8004 (
            .O(N__38635),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__8003 (
            .O(N__38632),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__8002 (
            .O(N__38625),
            .I(N__38622));
    InMux I__8001 (
            .O(N__38622),
            .I(N__38619));
    LocalMux I__8000 (
            .O(N__38619),
            .I(N__38616));
    Span4Mux_h I__7999 (
            .O(N__38616),
            .I(N__38613));
    Odrv4 I__7998 (
            .O(N__38613),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    InMux I__7997 (
            .O(N__38610),
            .I(N__38604));
    InMux I__7996 (
            .O(N__38609),
            .I(N__38604));
    LocalMux I__7995 (
            .O(N__38604),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    InMux I__7994 (
            .O(N__38601),
            .I(N__38598));
    LocalMux I__7993 (
            .O(N__38598),
            .I(N__38595));
    Odrv4 I__7992 (
            .O(N__38595),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__7991 (
            .O(N__38592),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__7990 (
            .O(N__38589),
            .I(N__38586));
    LocalMux I__7989 (
            .O(N__38586),
            .I(N__38583));
    Odrv4 I__7988 (
            .O(N__38583),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__7987 (
            .O(N__38580),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__7986 (
            .O(N__38577),
            .I(N__38574));
    LocalMux I__7985 (
            .O(N__38574),
            .I(N__38571));
    Odrv4 I__7984 (
            .O(N__38571),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__7983 (
            .O(N__38568),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__7982 (
            .O(N__38565),
            .I(N__38562));
    LocalMux I__7981 (
            .O(N__38562),
            .I(N__38559));
    Odrv4 I__7980 (
            .O(N__38559),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__7979 (
            .O(N__38556),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__7978 (
            .O(N__38553),
            .I(N__38550));
    LocalMux I__7977 (
            .O(N__38550),
            .I(N__38547));
    Odrv4 I__7976 (
            .O(N__38547),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__7975 (
            .O(N__38544),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__7974 (
            .O(N__38541),
            .I(N__38538));
    LocalMux I__7973 (
            .O(N__38538),
            .I(N__38535));
    Odrv4 I__7972 (
            .O(N__38535),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__7971 (
            .O(N__38532),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__7970 (
            .O(N__38529),
            .I(N__38525));
    InMux I__7969 (
            .O(N__38528),
            .I(N__38522));
    LocalMux I__7968 (
            .O(N__38525),
            .I(N__38515));
    LocalMux I__7967 (
            .O(N__38522),
            .I(N__38509));
    InMux I__7966 (
            .O(N__38521),
            .I(N__38500));
    InMux I__7965 (
            .O(N__38520),
            .I(N__38500));
    InMux I__7964 (
            .O(N__38519),
            .I(N__38500));
    InMux I__7963 (
            .O(N__38518),
            .I(N__38500));
    Span4Mux_h I__7962 (
            .O(N__38515),
            .I(N__38491));
    InMux I__7961 (
            .O(N__38514),
            .I(N__38484));
    InMux I__7960 (
            .O(N__38513),
            .I(N__38484));
    InMux I__7959 (
            .O(N__38512),
            .I(N__38484));
    Span4Mux_v I__7958 (
            .O(N__38509),
            .I(N__38479));
    LocalMux I__7957 (
            .O(N__38500),
            .I(N__38479));
    InMux I__7956 (
            .O(N__38499),
            .I(N__38468));
    InMux I__7955 (
            .O(N__38498),
            .I(N__38468));
    InMux I__7954 (
            .O(N__38497),
            .I(N__38468));
    InMux I__7953 (
            .O(N__38496),
            .I(N__38468));
    InMux I__7952 (
            .O(N__38495),
            .I(N__38468));
    InMux I__7951 (
            .O(N__38494),
            .I(N__38465));
    Odrv4 I__7950 (
            .O(N__38491),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__7949 (
            .O(N__38484),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__7948 (
            .O(N__38479),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__7947 (
            .O(N__38468),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__7946 (
            .O(N__38465),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__7945 (
            .O(N__38454),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__7944 (
            .O(N__38451),
            .I(N__38448));
    LocalMux I__7943 (
            .O(N__38448),
            .I(N__38445));
    Span4Mux_h I__7942 (
            .O(N__38445),
            .I(N__38442));
    Odrv4 I__7941 (
            .O(N__38442),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__7940 (
            .O(N__38439),
            .I(N__38436));
    LocalMux I__7939 (
            .O(N__38436),
            .I(N__38433));
    Span4Mux_h I__7938 (
            .O(N__38433),
            .I(N__38430));
    Odrv4 I__7937 (
            .O(N__38430),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    InMux I__7936 (
            .O(N__38427),
            .I(N__38424));
    LocalMux I__7935 (
            .O(N__38424),
            .I(N__38421));
    Odrv12 I__7934 (
            .O(N__38421),
            .I(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ));
    InMux I__7933 (
            .O(N__38418),
            .I(N__38415));
    LocalMux I__7932 (
            .O(N__38415),
            .I(N__38412));
    Span4Mux_h I__7931 (
            .O(N__38412),
            .I(N__38409));
    Odrv4 I__7930 (
            .O(N__38409),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__7929 (
            .O(N__38406),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__7928 (
            .O(N__38403),
            .I(N__38400));
    LocalMux I__7927 (
            .O(N__38400),
            .I(N__38397));
    Odrv4 I__7926 (
            .O(N__38397),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__7925 (
            .O(N__38394),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__7924 (
            .O(N__38391),
            .I(N__38388));
    LocalMux I__7923 (
            .O(N__38388),
            .I(N__38385));
    Odrv4 I__7922 (
            .O(N__38385),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__7921 (
            .O(N__38382),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__7920 (
            .O(N__38379),
            .I(N__38376));
    LocalMux I__7919 (
            .O(N__38376),
            .I(N__38373));
    Odrv4 I__7918 (
            .O(N__38373),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__7917 (
            .O(N__38370),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__7916 (
            .O(N__38367),
            .I(N__38364));
    LocalMux I__7915 (
            .O(N__38364),
            .I(N__38361));
    Odrv4 I__7914 (
            .O(N__38361),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__7913 (
            .O(N__38358),
            .I(bfn_15_15_0_));
    CascadeMux I__7912 (
            .O(N__38355),
            .I(N__38352));
    InMux I__7911 (
            .O(N__38352),
            .I(N__38349));
    LocalMux I__7910 (
            .O(N__38349),
            .I(N__38346));
    Span4Mux_v I__7909 (
            .O(N__38346),
            .I(N__38343));
    Odrv4 I__7908 (
            .O(N__38343),
            .I(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ));
    InMux I__7907 (
            .O(N__38340),
            .I(N__38337));
    LocalMux I__7906 (
            .O(N__38337),
            .I(N__38334));
    Span4Mux_v I__7905 (
            .O(N__38334),
            .I(N__38331));
    Odrv4 I__7904 (
            .O(N__38331),
            .I(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ));
    InMux I__7903 (
            .O(N__38328),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    CascadeMux I__7902 (
            .O(N__38325),
            .I(N__38322));
    InMux I__7901 (
            .O(N__38322),
            .I(N__38319));
    LocalMux I__7900 (
            .O(N__38319),
            .I(N__38316));
    Odrv12 I__7899 (
            .O(N__38316),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    InMux I__7898 (
            .O(N__38313),
            .I(N__38310));
    LocalMux I__7897 (
            .O(N__38310),
            .I(N__38307));
    Span4Mux_v I__7896 (
            .O(N__38307),
            .I(N__38304));
    Odrv4 I__7895 (
            .O(N__38304),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    InMux I__7894 (
            .O(N__38301),
            .I(N__38298));
    LocalMux I__7893 (
            .O(N__38298),
            .I(N__38295));
    Span4Mux_v I__7892 (
            .O(N__38295),
            .I(N__38292));
    Odrv4 I__7891 (
            .O(N__38292),
            .I(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ));
    InMux I__7890 (
            .O(N__38289),
            .I(N__38286));
    LocalMux I__7889 (
            .O(N__38286),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    InMux I__7888 (
            .O(N__38283),
            .I(N__38271));
    InMux I__7887 (
            .O(N__38282),
            .I(N__38267));
    InMux I__7886 (
            .O(N__38281),
            .I(N__38260));
    InMux I__7885 (
            .O(N__38280),
            .I(N__38260));
    InMux I__7884 (
            .O(N__38279),
            .I(N__38260));
    InMux I__7883 (
            .O(N__38278),
            .I(N__38251));
    InMux I__7882 (
            .O(N__38277),
            .I(N__38251));
    InMux I__7881 (
            .O(N__38276),
            .I(N__38251));
    InMux I__7880 (
            .O(N__38275),
            .I(N__38251));
    InMux I__7879 (
            .O(N__38274),
            .I(N__38240));
    LocalMux I__7878 (
            .O(N__38271),
            .I(N__38237));
    InMux I__7877 (
            .O(N__38270),
            .I(N__38233));
    LocalMux I__7876 (
            .O(N__38267),
            .I(N__38226));
    LocalMux I__7875 (
            .O(N__38260),
            .I(N__38226));
    LocalMux I__7874 (
            .O(N__38251),
            .I(N__38226));
    InMux I__7873 (
            .O(N__38250),
            .I(N__38223));
    InMux I__7872 (
            .O(N__38249),
            .I(N__38216));
    InMux I__7871 (
            .O(N__38248),
            .I(N__38216));
    InMux I__7870 (
            .O(N__38247),
            .I(N__38216));
    InMux I__7869 (
            .O(N__38246),
            .I(N__38207));
    InMux I__7868 (
            .O(N__38245),
            .I(N__38207));
    InMux I__7867 (
            .O(N__38244),
            .I(N__38207));
    InMux I__7866 (
            .O(N__38243),
            .I(N__38207));
    LocalMux I__7865 (
            .O(N__38240),
            .I(N__38204));
    Span4Mux_s2_h I__7864 (
            .O(N__38237),
            .I(N__38201));
    InMux I__7863 (
            .O(N__38236),
            .I(N__38195));
    LocalMux I__7862 (
            .O(N__38233),
            .I(N__38189));
    Span4Mux_v I__7861 (
            .O(N__38226),
            .I(N__38180));
    LocalMux I__7860 (
            .O(N__38223),
            .I(N__38180));
    LocalMux I__7859 (
            .O(N__38216),
            .I(N__38180));
    LocalMux I__7858 (
            .O(N__38207),
            .I(N__38180));
    Span12Mux_s2_h I__7857 (
            .O(N__38204),
            .I(N__38175));
    Sp12to4 I__7856 (
            .O(N__38201),
            .I(N__38175));
    InMux I__7855 (
            .O(N__38200),
            .I(N__38172));
    InMux I__7854 (
            .O(N__38199),
            .I(N__38167));
    InMux I__7853 (
            .O(N__38198),
            .I(N__38167));
    LocalMux I__7852 (
            .O(N__38195),
            .I(N__38164));
    CascadeMux I__7851 (
            .O(N__38194),
            .I(N__38158));
    CascadeMux I__7850 (
            .O(N__38193),
            .I(N__38154));
    CascadeMux I__7849 (
            .O(N__38192),
            .I(N__38150));
    Span12Mux_s6_h I__7848 (
            .O(N__38189),
            .I(N__38135));
    Span4Mux_v I__7847 (
            .O(N__38180),
            .I(N__38132));
    Span12Mux_v I__7846 (
            .O(N__38175),
            .I(N__38125));
    LocalMux I__7845 (
            .O(N__38172),
            .I(N__38125));
    LocalMux I__7844 (
            .O(N__38167),
            .I(N__38125));
    Span12Mux_s11_h I__7843 (
            .O(N__38164),
            .I(N__38122));
    InMux I__7842 (
            .O(N__38163),
            .I(N__38117));
    InMux I__7841 (
            .O(N__38162),
            .I(N__38117));
    InMux I__7840 (
            .O(N__38161),
            .I(N__38102));
    InMux I__7839 (
            .O(N__38158),
            .I(N__38102));
    InMux I__7838 (
            .O(N__38157),
            .I(N__38102));
    InMux I__7837 (
            .O(N__38154),
            .I(N__38102));
    InMux I__7836 (
            .O(N__38153),
            .I(N__38102));
    InMux I__7835 (
            .O(N__38150),
            .I(N__38102));
    InMux I__7834 (
            .O(N__38149),
            .I(N__38102));
    CascadeMux I__7833 (
            .O(N__38148),
            .I(N__38099));
    CascadeMux I__7832 (
            .O(N__38147),
            .I(N__38095));
    CascadeMux I__7831 (
            .O(N__38146),
            .I(N__38091));
    CascadeMux I__7830 (
            .O(N__38145),
            .I(N__38087));
    CascadeMux I__7829 (
            .O(N__38144),
            .I(N__38083));
    CascadeMux I__7828 (
            .O(N__38143),
            .I(N__38079));
    CascadeMux I__7827 (
            .O(N__38142),
            .I(N__38075));
    CascadeMux I__7826 (
            .O(N__38141),
            .I(N__38071));
    CascadeMux I__7825 (
            .O(N__38140),
            .I(N__38066));
    CascadeMux I__7824 (
            .O(N__38139),
            .I(N__38062));
    CascadeMux I__7823 (
            .O(N__38138),
            .I(N__38058));
    Span12Mux_v I__7822 (
            .O(N__38135),
            .I(N__38054));
    Sp12to4 I__7821 (
            .O(N__38132),
            .I(N__38051));
    Span12Mux_v I__7820 (
            .O(N__38125),
            .I(N__38048));
    Span12Mux_v I__7819 (
            .O(N__38122),
            .I(N__38043));
    LocalMux I__7818 (
            .O(N__38117),
            .I(N__38043));
    LocalMux I__7817 (
            .O(N__38102),
            .I(N__38040));
    InMux I__7816 (
            .O(N__38099),
            .I(N__38023));
    InMux I__7815 (
            .O(N__38098),
            .I(N__38023));
    InMux I__7814 (
            .O(N__38095),
            .I(N__38023));
    InMux I__7813 (
            .O(N__38094),
            .I(N__38023));
    InMux I__7812 (
            .O(N__38091),
            .I(N__38023));
    InMux I__7811 (
            .O(N__38090),
            .I(N__38023));
    InMux I__7810 (
            .O(N__38087),
            .I(N__38023));
    InMux I__7809 (
            .O(N__38086),
            .I(N__38023));
    InMux I__7808 (
            .O(N__38083),
            .I(N__38006));
    InMux I__7807 (
            .O(N__38082),
            .I(N__38006));
    InMux I__7806 (
            .O(N__38079),
            .I(N__38006));
    InMux I__7805 (
            .O(N__38078),
            .I(N__38006));
    InMux I__7804 (
            .O(N__38075),
            .I(N__38006));
    InMux I__7803 (
            .O(N__38074),
            .I(N__38006));
    InMux I__7802 (
            .O(N__38071),
            .I(N__38006));
    InMux I__7801 (
            .O(N__38070),
            .I(N__38006));
    InMux I__7800 (
            .O(N__38069),
            .I(N__37991));
    InMux I__7799 (
            .O(N__38066),
            .I(N__37991));
    InMux I__7798 (
            .O(N__38065),
            .I(N__37991));
    InMux I__7797 (
            .O(N__38062),
            .I(N__37991));
    InMux I__7796 (
            .O(N__38061),
            .I(N__37991));
    InMux I__7795 (
            .O(N__38058),
            .I(N__37991));
    InMux I__7794 (
            .O(N__38057),
            .I(N__37991));
    Span12Mux_v I__7793 (
            .O(N__38054),
            .I(N__37986));
    Span12Mux_s6_h I__7792 (
            .O(N__38051),
            .I(N__37986));
    Span12Mux_h I__7791 (
            .O(N__38048),
            .I(N__37981));
    Span12Mux_v I__7790 (
            .O(N__38043),
            .I(N__37981));
    Span12Mux_v I__7789 (
            .O(N__38040),
            .I(N__37972));
    LocalMux I__7788 (
            .O(N__38023),
            .I(N__37972));
    LocalMux I__7787 (
            .O(N__38006),
            .I(N__37972));
    LocalMux I__7786 (
            .O(N__37991),
            .I(N__37972));
    Odrv12 I__7785 (
            .O(N__37986),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__7784 (
            .O(N__37981),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__7783 (
            .O(N__37972),
            .I(CONSTANT_ONE_NET));
    InMux I__7782 (
            .O(N__37965),
            .I(N__37962));
    LocalMux I__7781 (
            .O(N__37962),
            .I(N__37959));
    Odrv4 I__7780 (
            .O(N__37959),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__7779 (
            .O(N__37956),
            .I(N__37953));
    InMux I__7778 (
            .O(N__37953),
            .I(N__37950));
    LocalMux I__7777 (
            .O(N__37950),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    InMux I__7776 (
            .O(N__37947),
            .I(N__37944));
    LocalMux I__7775 (
            .O(N__37944),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__7774 (
            .O(N__37941),
            .I(N__37938));
    LocalMux I__7773 (
            .O(N__37938),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    CascadeMux I__7772 (
            .O(N__37935),
            .I(N__37932));
    InMux I__7771 (
            .O(N__37932),
            .I(N__37929));
    LocalMux I__7770 (
            .O(N__37929),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__7769 (
            .O(N__37926),
            .I(N__37923));
    LocalMux I__7768 (
            .O(N__37923),
            .I(N__37919));
    InMux I__7767 (
            .O(N__37922),
            .I(N__37916));
    Sp12to4 I__7766 (
            .O(N__37919),
            .I(N__37910));
    LocalMux I__7765 (
            .O(N__37916),
            .I(N__37910));
    InMux I__7764 (
            .O(N__37915),
            .I(N__37907));
    Span12Mux_v I__7763 (
            .O(N__37910),
            .I(N__37904));
    LocalMux I__7762 (
            .O(N__37907),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    Odrv12 I__7761 (
            .O(N__37904),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    CascadeMux I__7760 (
            .O(N__37899),
            .I(N__37896));
    InMux I__7759 (
            .O(N__37896),
            .I(N__37892));
    InMux I__7758 (
            .O(N__37895),
            .I(N__37888));
    LocalMux I__7757 (
            .O(N__37892),
            .I(N__37885));
    CascadeMux I__7756 (
            .O(N__37891),
            .I(N__37882));
    LocalMux I__7755 (
            .O(N__37888),
            .I(N__37878));
    Span4Mux_v I__7754 (
            .O(N__37885),
            .I(N__37874));
    InMux I__7753 (
            .O(N__37882),
            .I(N__37869));
    InMux I__7752 (
            .O(N__37881),
            .I(N__37869));
    Span4Mux_v I__7751 (
            .O(N__37878),
            .I(N__37866));
    InMux I__7750 (
            .O(N__37877),
            .I(N__37863));
    Span4Mux_h I__7749 (
            .O(N__37874),
            .I(N__37860));
    LocalMux I__7748 (
            .O(N__37869),
            .I(N__37855));
    Span4Mux_h I__7747 (
            .O(N__37866),
            .I(N__37855));
    LocalMux I__7746 (
            .O(N__37863),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__7745 (
            .O(N__37860),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__7744 (
            .O(N__37855),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__7743 (
            .O(N__37848),
            .I(N__37845));
    LocalMux I__7742 (
            .O(N__37845),
            .I(N__37842));
    Span4Mux_h I__7741 (
            .O(N__37842),
            .I(N__37839));
    Span4Mux_v I__7740 (
            .O(N__37839),
            .I(N__37836));
    Odrv4 I__7739 (
            .O(N__37836),
            .I(\current_shift_inst.PI_CTRL.integrator_i_11 ));
    InMux I__7738 (
            .O(N__37833),
            .I(N__37829));
    InMux I__7737 (
            .O(N__37832),
            .I(N__37826));
    LocalMux I__7736 (
            .O(N__37829),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    LocalMux I__7735 (
            .O(N__37826),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__7734 (
            .O(N__37821),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__7733 (
            .O(N__37818),
            .I(N__37814));
    InMux I__7732 (
            .O(N__37817),
            .I(N__37811));
    LocalMux I__7731 (
            .O(N__37814),
            .I(N__37808));
    LocalMux I__7730 (
            .O(N__37811),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__7729 (
            .O(N__37808),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__7728 (
            .O(N__37803),
            .I(bfn_14_24_0_));
    InMux I__7727 (
            .O(N__37800),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__7726 (
            .O(N__37797),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__7725 (
            .O(N__37794),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__7724 (
            .O(N__37791),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__7723 (
            .O(N__37788),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__7722 (
            .O(N__37785),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__7721 (
            .O(N__37782),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__7720 (
            .O(N__37779),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__7719 (
            .O(N__37776),
            .I(bfn_14_23_0_));
    InMux I__7718 (
            .O(N__37773),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__7717 (
            .O(N__37770),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__7716 (
            .O(N__37767),
            .I(N__37763));
    InMux I__7715 (
            .O(N__37766),
            .I(N__37760));
    LocalMux I__7714 (
            .O(N__37763),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    LocalMux I__7713 (
            .O(N__37760),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__7712 (
            .O(N__37755),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__7711 (
            .O(N__37752),
            .I(N__37748));
    InMux I__7710 (
            .O(N__37751),
            .I(N__37745));
    LocalMux I__7709 (
            .O(N__37748),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    LocalMux I__7708 (
            .O(N__37745),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__7707 (
            .O(N__37740),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__7706 (
            .O(N__37737),
            .I(N__37733));
    InMux I__7705 (
            .O(N__37736),
            .I(N__37730));
    LocalMux I__7704 (
            .O(N__37733),
            .I(N__37727));
    LocalMux I__7703 (
            .O(N__37730),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__7702 (
            .O(N__37727),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__7701 (
            .O(N__37722),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__7700 (
            .O(N__37719),
            .I(N__37716));
    LocalMux I__7699 (
            .O(N__37716),
            .I(N__37712));
    InMux I__7698 (
            .O(N__37715),
            .I(N__37709));
    Span4Mux_h I__7697 (
            .O(N__37712),
            .I(N__37706));
    LocalMux I__7696 (
            .O(N__37709),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__7695 (
            .O(N__37706),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__7694 (
            .O(N__37701),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__7693 (
            .O(N__37698),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__7692 (
            .O(N__37695),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__7691 (
            .O(N__37692),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__7690 (
            .O(N__37689),
            .I(bfn_14_22_0_));
    InMux I__7689 (
            .O(N__37686),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__7688 (
            .O(N__37683),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__7687 (
            .O(N__37680),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__7686 (
            .O(N__37677),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__7685 (
            .O(N__37674),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    CascadeMux I__7684 (
            .O(N__37671),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__7683 (
            .O(N__37668),
            .I(N__37662));
    InMux I__7682 (
            .O(N__37667),
            .I(N__37662));
    LocalMux I__7681 (
            .O(N__37662),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__7680 (
            .O(N__37659),
            .I(N__37656));
    InMux I__7679 (
            .O(N__37656),
            .I(N__37649));
    InMux I__7678 (
            .O(N__37655),
            .I(N__37644));
    InMux I__7677 (
            .O(N__37654),
            .I(N__37644));
    InMux I__7676 (
            .O(N__37653),
            .I(N__37639));
    InMux I__7675 (
            .O(N__37652),
            .I(N__37639));
    LocalMux I__7674 (
            .O(N__37649),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__7673 (
            .O(N__37644),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__7672 (
            .O(N__37639),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    CascadeMux I__7671 (
            .O(N__37632),
            .I(N__37627));
    InMux I__7670 (
            .O(N__37631),
            .I(N__37622));
    InMux I__7669 (
            .O(N__37630),
            .I(N__37613));
    InMux I__7668 (
            .O(N__37627),
            .I(N__37613));
    InMux I__7667 (
            .O(N__37626),
            .I(N__37613));
    InMux I__7666 (
            .O(N__37625),
            .I(N__37613));
    LocalMux I__7665 (
            .O(N__37622),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__7664 (
            .O(N__37613),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__7663 (
            .O(N__37608),
            .I(N__37604));
    InMux I__7662 (
            .O(N__37607),
            .I(N__37601));
    LocalMux I__7661 (
            .O(N__37604),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    LocalMux I__7660 (
            .O(N__37601),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    InMux I__7659 (
            .O(N__37596),
            .I(N__37593));
    LocalMux I__7658 (
            .O(N__37593),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    InMux I__7657 (
            .O(N__37590),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__7656 (
            .O(N__37587),
            .I(N__37584));
    InMux I__7655 (
            .O(N__37584),
            .I(N__37581));
    LocalMux I__7654 (
            .O(N__37581),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28 ));
    InMux I__7653 (
            .O(N__37578),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__7652 (
            .O(N__37575),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__7651 (
            .O(N__37572),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__7650 (
            .O(N__37569),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__7649 (
            .O(N__37566),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__7648 (
            .O(N__37563),
            .I(N__37560));
    LocalMux I__7647 (
            .O(N__37560),
            .I(N__37556));
    InMux I__7646 (
            .O(N__37559),
            .I(N__37553));
    Span4Mux_h I__7645 (
            .O(N__37556),
            .I(N__37550));
    LocalMux I__7644 (
            .O(N__37553),
            .I(N__37547));
    Sp12to4 I__7643 (
            .O(N__37550),
            .I(N__37540));
    Sp12to4 I__7642 (
            .O(N__37547),
            .I(N__37540));
    InMux I__7641 (
            .O(N__37546),
            .I(N__37535));
    InMux I__7640 (
            .O(N__37545),
            .I(N__37535));
    Span12Mux_v I__7639 (
            .O(N__37540),
            .I(N__37532));
    LocalMux I__7638 (
            .O(N__37535),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv12 I__7637 (
            .O(N__37532),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__7636 (
            .O(N__37527),
            .I(N__37524));
    LocalMux I__7635 (
            .O(N__37524),
            .I(N__37520));
    InMux I__7634 (
            .O(N__37523),
            .I(N__37517));
    Span4Mux_v I__7633 (
            .O(N__37520),
            .I(N__37514));
    LocalMux I__7632 (
            .O(N__37517),
            .I(N__37511));
    Span4Mux_v I__7631 (
            .O(N__37514),
            .I(N__37508));
    Span12Mux_v I__7630 (
            .O(N__37511),
            .I(N__37504));
    Span4Mux_v I__7629 (
            .O(N__37508),
            .I(N__37501));
    InMux I__7628 (
            .O(N__37507),
            .I(N__37498));
    Odrv12 I__7627 (
            .O(N__37504),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__7626 (
            .O(N__37501),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    LocalMux I__7625 (
            .O(N__37498),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    CascadeMux I__7624 (
            .O(N__37491),
            .I(N__37488));
    InMux I__7623 (
            .O(N__37488),
            .I(N__37485));
    LocalMux I__7622 (
            .O(N__37485),
            .I(N__37479));
    InMux I__7621 (
            .O(N__37484),
            .I(N__37476));
    InMux I__7620 (
            .O(N__37483),
            .I(N__37473));
    InMux I__7619 (
            .O(N__37482),
            .I(N__37470));
    Span4Mux_h I__7618 (
            .O(N__37479),
            .I(N__37467));
    LocalMux I__7617 (
            .O(N__37476),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__7616 (
            .O(N__37473),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__7615 (
            .O(N__37470),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__7614 (
            .O(N__37467),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__7613 (
            .O(N__37458),
            .I(N__37453));
    InMux I__7612 (
            .O(N__37457),
            .I(N__37450));
    InMux I__7611 (
            .O(N__37456),
            .I(N__37447));
    LocalMux I__7610 (
            .O(N__37453),
            .I(N__37444));
    LocalMux I__7609 (
            .O(N__37450),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__7608 (
            .O(N__37447),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__7607 (
            .O(N__37444),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    CascadeMux I__7606 (
            .O(N__37437),
            .I(N__37434));
    InMux I__7605 (
            .O(N__37434),
            .I(N__37431));
    LocalMux I__7604 (
            .O(N__37431),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    InMux I__7603 (
            .O(N__37428),
            .I(N__37424));
    InMux I__7602 (
            .O(N__37427),
            .I(N__37421));
    LocalMux I__7601 (
            .O(N__37424),
            .I(N__37418));
    LocalMux I__7600 (
            .O(N__37421),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__7599 (
            .O(N__37418),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__7598 (
            .O(N__37413),
            .I(N__37409));
    InMux I__7597 (
            .O(N__37412),
            .I(N__37406));
    LocalMux I__7596 (
            .O(N__37409),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    LocalMux I__7595 (
            .O(N__37406),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__7594 (
            .O(N__37401),
            .I(N__37398));
    LocalMux I__7593 (
            .O(N__37398),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df24 ));
    CascadeMux I__7592 (
            .O(N__37395),
            .I(N__37392));
    InMux I__7591 (
            .O(N__37392),
            .I(N__37389));
    LocalMux I__7590 (
            .O(N__37389),
            .I(N__37386));
    Span4Mux_v I__7589 (
            .O(N__37386),
            .I(N__37383));
    Odrv4 I__7588 (
            .O(N__37383),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    InMux I__7587 (
            .O(N__37380),
            .I(N__37377));
    LocalMux I__7586 (
            .O(N__37377),
            .I(N__37374));
    Odrv4 I__7585 (
            .O(N__37374),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    InMux I__7584 (
            .O(N__37371),
            .I(N__37368));
    LocalMux I__7583 (
            .O(N__37368),
            .I(N__37365));
    Span4Mux_h I__7582 (
            .O(N__37365),
            .I(N__37362));
    Odrv4 I__7581 (
            .O(N__37362),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    InMux I__7580 (
            .O(N__37359),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__7579 (
            .O(N__37356),
            .I(N__37352));
    InMux I__7578 (
            .O(N__37355),
            .I(N__37349));
    LocalMux I__7577 (
            .O(N__37352),
            .I(N__37346));
    LocalMux I__7576 (
            .O(N__37349),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__7575 (
            .O(N__37346),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__7574 (
            .O(N__37341),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__7573 (
            .O(N__37338),
            .I(N__37334));
    InMux I__7572 (
            .O(N__37337),
            .I(N__37331));
    LocalMux I__7571 (
            .O(N__37334),
            .I(N__37328));
    LocalMux I__7570 (
            .O(N__37331),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__7569 (
            .O(N__37328),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__7568 (
            .O(N__37323),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__7567 (
            .O(N__37320),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__7566 (
            .O(N__37317),
            .I(bfn_14_17_0_));
    InMux I__7565 (
            .O(N__37314),
            .I(N__37311));
    LocalMux I__7564 (
            .O(N__37311),
            .I(N__37308));
    Span4Mux_v I__7563 (
            .O(N__37308),
            .I(N__37304));
    InMux I__7562 (
            .O(N__37307),
            .I(N__37301));
    Span4Mux_v I__7561 (
            .O(N__37304),
            .I(N__37298));
    LocalMux I__7560 (
            .O(N__37301),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv4 I__7559 (
            .O(N__37298),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__7558 (
            .O(N__37293),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__7557 (
            .O(N__37290),
            .I(N__37287));
    LocalMux I__7556 (
            .O(N__37287),
            .I(N__37284));
    Span4Mux_h I__7555 (
            .O(N__37284),
            .I(N__37280));
    InMux I__7554 (
            .O(N__37283),
            .I(N__37277));
    Span4Mux_v I__7553 (
            .O(N__37280),
            .I(N__37274));
    LocalMux I__7552 (
            .O(N__37277),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__7551 (
            .O(N__37274),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__7550 (
            .O(N__37269),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__7549 (
            .O(N__37266),
            .I(N__37263));
    LocalMux I__7548 (
            .O(N__37263),
            .I(N__37260));
    Span4Mux_h I__7547 (
            .O(N__37260),
            .I(N__37256));
    InMux I__7546 (
            .O(N__37259),
            .I(N__37253));
    Span4Mux_v I__7545 (
            .O(N__37256),
            .I(N__37250));
    LocalMux I__7544 (
            .O(N__37253),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__7543 (
            .O(N__37250),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__7542 (
            .O(N__37245),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__7541 (
            .O(N__37242),
            .I(N__37239));
    LocalMux I__7540 (
            .O(N__37239),
            .I(N__37236));
    Span4Mux_h I__7539 (
            .O(N__37236),
            .I(N__37232));
    InMux I__7538 (
            .O(N__37235),
            .I(N__37229));
    Span4Mux_v I__7537 (
            .O(N__37232),
            .I(N__37226));
    LocalMux I__7536 (
            .O(N__37229),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__7535 (
            .O(N__37226),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__7534 (
            .O(N__37221),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__7533 (
            .O(N__37218),
            .I(N__37214));
    InMux I__7532 (
            .O(N__37217),
            .I(N__37211));
    LocalMux I__7531 (
            .O(N__37214),
            .I(N__37208));
    LocalMux I__7530 (
            .O(N__37211),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__7529 (
            .O(N__37208),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__7528 (
            .O(N__37203),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__7527 (
            .O(N__37200),
            .I(N__37196));
    InMux I__7526 (
            .O(N__37199),
            .I(N__37193));
    LocalMux I__7525 (
            .O(N__37196),
            .I(N__37190));
    LocalMux I__7524 (
            .O(N__37193),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__7523 (
            .O(N__37190),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__7522 (
            .O(N__37185),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__7521 (
            .O(N__37182),
            .I(N__37178));
    InMux I__7520 (
            .O(N__37181),
            .I(N__37175));
    LocalMux I__7519 (
            .O(N__37178),
            .I(N__37172));
    LocalMux I__7518 (
            .O(N__37175),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__7517 (
            .O(N__37172),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__7516 (
            .O(N__37167),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__7515 (
            .O(N__37164),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__7514 (
            .O(N__37161),
            .I(bfn_14_16_0_));
    InMux I__7513 (
            .O(N__37158),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__7512 (
            .O(N__37155),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__7511 (
            .O(N__37152),
            .I(N__37148));
    InMux I__7510 (
            .O(N__37151),
            .I(N__37145));
    LocalMux I__7509 (
            .O(N__37148),
            .I(N__37142));
    LocalMux I__7508 (
            .O(N__37145),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__7507 (
            .O(N__37142),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__7506 (
            .O(N__37137),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__7505 (
            .O(N__37134),
            .I(N__37130));
    InMux I__7504 (
            .O(N__37133),
            .I(N__37127));
    LocalMux I__7503 (
            .O(N__37130),
            .I(N__37124));
    LocalMux I__7502 (
            .O(N__37127),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__7501 (
            .O(N__37124),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__7500 (
            .O(N__37119),
            .I(N__37115));
    InMux I__7499 (
            .O(N__37118),
            .I(N__37112));
    LocalMux I__7498 (
            .O(N__37115),
            .I(N__37109));
    LocalMux I__7497 (
            .O(N__37112),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__7496 (
            .O(N__37109),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__7495 (
            .O(N__37104),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__7494 (
            .O(N__37101),
            .I(N__37097));
    InMux I__7493 (
            .O(N__37100),
            .I(N__37094));
    LocalMux I__7492 (
            .O(N__37097),
            .I(N__37091));
    LocalMux I__7491 (
            .O(N__37094),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__7490 (
            .O(N__37091),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__7489 (
            .O(N__37086),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__7488 (
            .O(N__37083),
            .I(N__37079));
    InMux I__7487 (
            .O(N__37082),
            .I(N__37076));
    LocalMux I__7486 (
            .O(N__37079),
            .I(N__37073));
    LocalMux I__7485 (
            .O(N__37076),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__7484 (
            .O(N__37073),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__7483 (
            .O(N__37068),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__7482 (
            .O(N__37065),
            .I(N__37061));
    InMux I__7481 (
            .O(N__37064),
            .I(N__37058));
    LocalMux I__7480 (
            .O(N__37061),
            .I(N__37055));
    LocalMux I__7479 (
            .O(N__37058),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__7478 (
            .O(N__37055),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__7477 (
            .O(N__37050),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__7476 (
            .O(N__37047),
            .I(N__37043));
    InMux I__7475 (
            .O(N__37046),
            .I(N__37040));
    LocalMux I__7474 (
            .O(N__37043),
            .I(N__37037));
    LocalMux I__7473 (
            .O(N__37040),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__7472 (
            .O(N__37037),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__7471 (
            .O(N__37032),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__7470 (
            .O(N__37029),
            .I(N__37025));
    InMux I__7469 (
            .O(N__37028),
            .I(N__37022));
    LocalMux I__7468 (
            .O(N__37025),
            .I(N__37019));
    LocalMux I__7467 (
            .O(N__37022),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__7466 (
            .O(N__37019),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__7465 (
            .O(N__37014),
            .I(bfn_14_15_0_));
    InMux I__7464 (
            .O(N__37011),
            .I(N__37008));
    LocalMux I__7463 (
            .O(N__37008),
            .I(N__37004));
    InMux I__7462 (
            .O(N__37007),
            .I(N__37001));
    Span4Mux_v I__7461 (
            .O(N__37004),
            .I(N__36998));
    LocalMux I__7460 (
            .O(N__37001),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__7459 (
            .O(N__36998),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__7458 (
            .O(N__36993),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__7457 (
            .O(N__36990),
            .I(N__36986));
    InMux I__7456 (
            .O(N__36989),
            .I(N__36983));
    LocalMux I__7455 (
            .O(N__36986),
            .I(N__36980));
    LocalMux I__7454 (
            .O(N__36983),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__7453 (
            .O(N__36980),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__7452 (
            .O(N__36975),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__7451 (
            .O(N__36972),
            .I(N__36968));
    InMux I__7450 (
            .O(N__36971),
            .I(N__36965));
    LocalMux I__7449 (
            .O(N__36968),
            .I(N__36962));
    LocalMux I__7448 (
            .O(N__36965),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__7447 (
            .O(N__36962),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__7446 (
            .O(N__36957),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__7445 (
            .O(N__36954),
            .I(N__36951));
    LocalMux I__7444 (
            .O(N__36951),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__7443 (
            .O(N__36948),
            .I(N__36945));
    LocalMux I__7442 (
            .O(N__36945),
            .I(N__36942));
    Odrv4 I__7441 (
            .O(N__36942),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__7440 (
            .O(N__36939),
            .I(N__36936));
    LocalMux I__7439 (
            .O(N__36936),
            .I(N__36933));
    Odrv4 I__7438 (
            .O(N__36933),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__7437 (
            .O(N__36930),
            .I(N__36927));
    LocalMux I__7436 (
            .O(N__36927),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__7435 (
            .O(N__36924),
            .I(N__36921));
    LocalMux I__7434 (
            .O(N__36921),
            .I(\current_shift_inst.control_input_axb_10 ));
    CascadeMux I__7433 (
            .O(N__36918),
            .I(N__36915));
    InMux I__7432 (
            .O(N__36915),
            .I(N__36910));
    InMux I__7431 (
            .O(N__36914),
            .I(N__36907));
    InMux I__7430 (
            .O(N__36913),
            .I(N__36904));
    LocalMux I__7429 (
            .O(N__36910),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__7428 (
            .O(N__36907),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__7427 (
            .O(N__36904),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__7426 (
            .O(N__36897),
            .I(N__36894));
    InMux I__7425 (
            .O(N__36894),
            .I(N__36891));
    LocalMux I__7424 (
            .O(N__36891),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    InMux I__7423 (
            .O(N__36888),
            .I(N__36884));
    InMux I__7422 (
            .O(N__36887),
            .I(N__36881));
    LocalMux I__7421 (
            .O(N__36884),
            .I(N__36878));
    LocalMux I__7420 (
            .O(N__36881),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__7419 (
            .O(N__36878),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__7418 (
            .O(N__36873),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__7417 (
            .O(N__36870),
            .I(N__36867));
    InMux I__7416 (
            .O(N__36867),
            .I(N__36864));
    LocalMux I__7415 (
            .O(N__36864),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28 ));
    InMux I__7414 (
            .O(N__36861),
            .I(N__36857));
    InMux I__7413 (
            .O(N__36860),
            .I(N__36854));
    LocalMux I__7412 (
            .O(N__36857),
            .I(N__36851));
    LocalMux I__7411 (
            .O(N__36854),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__7410 (
            .O(N__36851),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__7409 (
            .O(N__36846),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    CascadeMux I__7408 (
            .O(N__36843),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    InMux I__7407 (
            .O(N__36840),
            .I(N__36837));
    LocalMux I__7406 (
            .O(N__36837),
            .I(N__36833));
    InMux I__7405 (
            .O(N__36836),
            .I(N__36830));
    Span4Mux_h I__7404 (
            .O(N__36833),
            .I(N__36827));
    LocalMux I__7403 (
            .O(N__36830),
            .I(N__36824));
    Span4Mux_h I__7402 (
            .O(N__36827),
            .I(N__36821));
    Span4Mux_h I__7401 (
            .O(N__36824),
            .I(N__36818));
    Odrv4 I__7400 (
            .O(N__36821),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv4 I__7399 (
            .O(N__36818),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__7398 (
            .O(N__36813),
            .I(N__36810));
    LocalMux I__7397 (
            .O(N__36810),
            .I(N__36807));
    Odrv4 I__7396 (
            .O(N__36807),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    InMux I__7395 (
            .O(N__36804),
            .I(N__36801));
    LocalMux I__7394 (
            .O(N__36801),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__7393 (
            .O(N__36798),
            .I(N__36795));
    LocalMux I__7392 (
            .O(N__36795),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__7391 (
            .O(N__36792),
            .I(N__36788));
    CascadeMux I__7390 (
            .O(N__36791),
            .I(N__36784));
    LocalMux I__7389 (
            .O(N__36788),
            .I(N__36781));
    InMux I__7388 (
            .O(N__36787),
            .I(N__36778));
    InMux I__7387 (
            .O(N__36784),
            .I(N__36775));
    Odrv4 I__7386 (
            .O(N__36781),
            .I(\current_shift_inst.N_1460_i ));
    LocalMux I__7385 (
            .O(N__36778),
            .I(\current_shift_inst.N_1460_i ));
    LocalMux I__7384 (
            .O(N__36775),
            .I(\current_shift_inst.N_1460_i ));
    InMux I__7383 (
            .O(N__36768),
            .I(N__36765));
    LocalMux I__7382 (
            .O(N__36765),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__7381 (
            .O(N__36762),
            .I(N__36759));
    LocalMux I__7380 (
            .O(N__36759),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__7379 (
            .O(N__36756),
            .I(N__36753));
    LocalMux I__7378 (
            .O(N__36753),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__7377 (
            .O(N__36750),
            .I(N__36747));
    LocalMux I__7376 (
            .O(N__36747),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__7375 (
            .O(N__36744),
            .I(N__36741));
    LocalMux I__7374 (
            .O(N__36741),
            .I(\current_shift_inst.control_input_axb_0 ));
    CascadeMux I__7373 (
            .O(N__36738),
            .I(N__36734));
    CascadeMux I__7372 (
            .O(N__36737),
            .I(N__36731));
    InMux I__7371 (
            .O(N__36734),
            .I(N__36725));
    InMux I__7370 (
            .O(N__36731),
            .I(N__36725));
    InMux I__7369 (
            .O(N__36730),
            .I(N__36722));
    LocalMux I__7368 (
            .O(N__36725),
            .I(N__36719));
    LocalMux I__7367 (
            .O(N__36722),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__7366 (
            .O(N__36719),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__7365 (
            .O(N__36714),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__7364 (
            .O(N__36711),
            .I(N__36704));
    InMux I__7363 (
            .O(N__36710),
            .I(N__36704));
    InMux I__7362 (
            .O(N__36709),
            .I(N__36701));
    LocalMux I__7361 (
            .O(N__36704),
            .I(N__36698));
    LocalMux I__7360 (
            .O(N__36701),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__7359 (
            .O(N__36698),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__7358 (
            .O(N__36693),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__7357 (
            .O(N__36690),
            .I(N__36686));
    InMux I__7356 (
            .O(N__36689),
            .I(N__36683));
    LocalMux I__7355 (
            .O(N__36686),
            .I(N__36680));
    LocalMux I__7354 (
            .O(N__36683),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__7353 (
            .O(N__36680),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__7352 (
            .O(N__36675),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__7351 (
            .O(N__36672),
            .I(N__36658));
    InMux I__7350 (
            .O(N__36671),
            .I(N__36658));
    InMux I__7349 (
            .O(N__36670),
            .I(N__36637));
    InMux I__7348 (
            .O(N__36669),
            .I(N__36637));
    InMux I__7347 (
            .O(N__36668),
            .I(N__36637));
    InMux I__7346 (
            .O(N__36667),
            .I(N__36637));
    InMux I__7345 (
            .O(N__36666),
            .I(N__36620));
    InMux I__7344 (
            .O(N__36665),
            .I(N__36620));
    InMux I__7343 (
            .O(N__36664),
            .I(N__36620));
    InMux I__7342 (
            .O(N__36663),
            .I(N__36620));
    LocalMux I__7341 (
            .O(N__36658),
            .I(N__36617));
    InMux I__7340 (
            .O(N__36657),
            .I(N__36608));
    InMux I__7339 (
            .O(N__36656),
            .I(N__36608));
    InMux I__7338 (
            .O(N__36655),
            .I(N__36608));
    InMux I__7337 (
            .O(N__36654),
            .I(N__36608));
    InMux I__7336 (
            .O(N__36653),
            .I(N__36599));
    InMux I__7335 (
            .O(N__36652),
            .I(N__36599));
    InMux I__7334 (
            .O(N__36651),
            .I(N__36599));
    InMux I__7333 (
            .O(N__36650),
            .I(N__36599));
    InMux I__7332 (
            .O(N__36649),
            .I(N__36590));
    InMux I__7331 (
            .O(N__36648),
            .I(N__36590));
    InMux I__7330 (
            .O(N__36647),
            .I(N__36590));
    InMux I__7329 (
            .O(N__36646),
            .I(N__36590));
    LocalMux I__7328 (
            .O(N__36637),
            .I(N__36587));
    InMux I__7327 (
            .O(N__36636),
            .I(N__36578));
    InMux I__7326 (
            .O(N__36635),
            .I(N__36578));
    InMux I__7325 (
            .O(N__36634),
            .I(N__36578));
    InMux I__7324 (
            .O(N__36633),
            .I(N__36578));
    InMux I__7323 (
            .O(N__36632),
            .I(N__36569));
    InMux I__7322 (
            .O(N__36631),
            .I(N__36569));
    InMux I__7321 (
            .O(N__36630),
            .I(N__36569));
    InMux I__7320 (
            .O(N__36629),
            .I(N__36569));
    LocalMux I__7319 (
            .O(N__36620),
            .I(N__36558));
    Span4Mux_h I__7318 (
            .O(N__36617),
            .I(N__36558));
    LocalMux I__7317 (
            .O(N__36608),
            .I(N__36558));
    LocalMux I__7316 (
            .O(N__36599),
            .I(N__36558));
    LocalMux I__7315 (
            .O(N__36590),
            .I(N__36558));
    Odrv4 I__7314 (
            .O(N__36587),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__7313 (
            .O(N__36578),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__7312 (
            .O(N__36569),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__7311 (
            .O(N__36558),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__7310 (
            .O(N__36549),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CascadeMux I__7309 (
            .O(N__36546),
            .I(N__36543));
    InMux I__7308 (
            .O(N__36543),
            .I(N__36539));
    InMux I__7307 (
            .O(N__36542),
            .I(N__36536));
    LocalMux I__7306 (
            .O(N__36539),
            .I(N__36533));
    LocalMux I__7305 (
            .O(N__36536),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__7304 (
            .O(N__36533),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__7303 (
            .O(N__36528),
            .I(N__36525));
    LocalMux I__7302 (
            .O(N__36525),
            .I(N__36520));
    CEMux I__7301 (
            .O(N__36524),
            .I(N__36517));
    CEMux I__7300 (
            .O(N__36523),
            .I(N__36513));
    Span4Mux_v I__7299 (
            .O(N__36520),
            .I(N__36508));
    LocalMux I__7298 (
            .O(N__36517),
            .I(N__36508));
    CEMux I__7297 (
            .O(N__36516),
            .I(N__36505));
    LocalMux I__7296 (
            .O(N__36513),
            .I(N__36502));
    Span4Mux_v I__7295 (
            .O(N__36508),
            .I(N__36497));
    LocalMux I__7294 (
            .O(N__36505),
            .I(N__36497));
    Span4Mux_v I__7293 (
            .O(N__36502),
            .I(N__36494));
    Span4Mux_v I__7292 (
            .O(N__36497),
            .I(N__36489));
    Span4Mux_s1_v I__7291 (
            .O(N__36494),
            .I(N__36489));
    Odrv4 I__7290 (
            .O(N__36489),
            .I(\current_shift_inst.timer_s1.N_167_i ));
    CascadeMux I__7289 (
            .O(N__36486),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_ ));
    CascadeMux I__7288 (
            .O(N__36483),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    CascadeMux I__7287 (
            .O(N__36480),
            .I(N__36477));
    InMux I__7286 (
            .O(N__36477),
            .I(N__36474));
    LocalMux I__7285 (
            .O(N__36474),
            .I(N__36470));
    InMux I__7284 (
            .O(N__36473),
            .I(N__36466));
    Span4Mux_h I__7283 (
            .O(N__36470),
            .I(N__36463));
    InMux I__7282 (
            .O(N__36469),
            .I(N__36460));
    LocalMux I__7281 (
            .O(N__36466),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__7280 (
            .O(N__36463),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    LocalMux I__7279 (
            .O(N__36460),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__7278 (
            .O(N__36453),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__7277 (
            .O(N__36450),
            .I(N__36444));
    InMux I__7276 (
            .O(N__36449),
            .I(N__36444));
    LocalMux I__7275 (
            .O(N__36444),
            .I(N__36440));
    InMux I__7274 (
            .O(N__36443),
            .I(N__36437));
    Span4Mux_v I__7273 (
            .O(N__36440),
            .I(N__36434));
    LocalMux I__7272 (
            .O(N__36437),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__7271 (
            .O(N__36434),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__7270 (
            .O(N__36429),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__7269 (
            .O(N__36426),
            .I(N__36419));
    InMux I__7268 (
            .O(N__36425),
            .I(N__36419));
    InMux I__7267 (
            .O(N__36424),
            .I(N__36416));
    LocalMux I__7266 (
            .O(N__36419),
            .I(N__36413));
    LocalMux I__7265 (
            .O(N__36416),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__7264 (
            .O(N__36413),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__7263 (
            .O(N__36408),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__7262 (
            .O(N__36405),
            .I(N__36401));
    CascadeMux I__7261 (
            .O(N__36404),
            .I(N__36398));
    InMux I__7260 (
            .O(N__36401),
            .I(N__36393));
    InMux I__7259 (
            .O(N__36398),
            .I(N__36393));
    LocalMux I__7258 (
            .O(N__36393),
            .I(N__36389));
    InMux I__7257 (
            .O(N__36392),
            .I(N__36386));
    Span4Mux_h I__7256 (
            .O(N__36389),
            .I(N__36383));
    LocalMux I__7255 (
            .O(N__36386),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__7254 (
            .O(N__36383),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__7253 (
            .O(N__36378),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__7252 (
            .O(N__36375),
            .I(N__36371));
    CascadeMux I__7251 (
            .O(N__36374),
            .I(N__36368));
    InMux I__7250 (
            .O(N__36371),
            .I(N__36362));
    InMux I__7249 (
            .O(N__36368),
            .I(N__36362));
    InMux I__7248 (
            .O(N__36367),
            .I(N__36359));
    LocalMux I__7247 (
            .O(N__36362),
            .I(N__36356));
    LocalMux I__7246 (
            .O(N__36359),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__7245 (
            .O(N__36356),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__7244 (
            .O(N__36351),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__7243 (
            .O(N__36348),
            .I(N__36341));
    InMux I__7242 (
            .O(N__36347),
            .I(N__36341));
    InMux I__7241 (
            .O(N__36346),
            .I(N__36338));
    LocalMux I__7240 (
            .O(N__36341),
            .I(N__36335));
    LocalMux I__7239 (
            .O(N__36338),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__7238 (
            .O(N__36335),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__7237 (
            .O(N__36330),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__7236 (
            .O(N__36327),
            .I(N__36323));
    InMux I__7235 (
            .O(N__36326),
            .I(N__36320));
    InMux I__7234 (
            .O(N__36323),
            .I(N__36316));
    LocalMux I__7233 (
            .O(N__36320),
            .I(N__36313));
    InMux I__7232 (
            .O(N__36319),
            .I(N__36310));
    LocalMux I__7231 (
            .O(N__36316),
            .I(N__36305));
    Span4Mux_h I__7230 (
            .O(N__36313),
            .I(N__36305));
    LocalMux I__7229 (
            .O(N__36310),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__7228 (
            .O(N__36305),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__7227 (
            .O(N__36300),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__7226 (
            .O(N__36297),
            .I(N__36294));
    LocalMux I__7225 (
            .O(N__36294),
            .I(N__36289));
    CascadeMux I__7224 (
            .O(N__36293),
            .I(N__36286));
    InMux I__7223 (
            .O(N__36292),
            .I(N__36283));
    Span4Mux_h I__7222 (
            .O(N__36289),
            .I(N__36280));
    InMux I__7221 (
            .O(N__36286),
            .I(N__36277));
    LocalMux I__7220 (
            .O(N__36283),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__7219 (
            .O(N__36280),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    LocalMux I__7218 (
            .O(N__36277),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__7217 (
            .O(N__36270),
            .I(bfn_14_8_0_));
    CascadeMux I__7216 (
            .O(N__36267),
            .I(N__36264));
    InMux I__7215 (
            .O(N__36264),
            .I(N__36261));
    LocalMux I__7214 (
            .O(N__36261),
            .I(N__36257));
    InMux I__7213 (
            .O(N__36260),
            .I(N__36253));
    Span4Mux_h I__7212 (
            .O(N__36257),
            .I(N__36250));
    InMux I__7211 (
            .O(N__36256),
            .I(N__36247));
    LocalMux I__7210 (
            .O(N__36253),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__7209 (
            .O(N__36250),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    LocalMux I__7208 (
            .O(N__36247),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__7207 (
            .O(N__36240),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__7206 (
            .O(N__36237),
            .I(N__36234));
    InMux I__7205 (
            .O(N__36234),
            .I(N__36231));
    LocalMux I__7204 (
            .O(N__36231),
            .I(N__36227));
    InMux I__7203 (
            .O(N__36230),
            .I(N__36223));
    Span4Mux_h I__7202 (
            .O(N__36227),
            .I(N__36220));
    InMux I__7201 (
            .O(N__36226),
            .I(N__36217));
    LocalMux I__7200 (
            .O(N__36223),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__7199 (
            .O(N__36220),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    LocalMux I__7198 (
            .O(N__36217),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__7197 (
            .O(N__36210),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__7196 (
            .O(N__36207),
            .I(N__36201));
    InMux I__7195 (
            .O(N__36206),
            .I(N__36201));
    LocalMux I__7194 (
            .O(N__36201),
            .I(N__36197));
    InMux I__7193 (
            .O(N__36200),
            .I(N__36194));
    Span4Mux_v I__7192 (
            .O(N__36197),
            .I(N__36191));
    LocalMux I__7191 (
            .O(N__36194),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__7190 (
            .O(N__36191),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__7189 (
            .O(N__36186),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__7188 (
            .O(N__36183),
            .I(N__36176));
    InMux I__7187 (
            .O(N__36182),
            .I(N__36176));
    InMux I__7186 (
            .O(N__36181),
            .I(N__36173));
    LocalMux I__7185 (
            .O(N__36176),
            .I(N__36170));
    LocalMux I__7184 (
            .O(N__36173),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__7183 (
            .O(N__36170),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__7182 (
            .O(N__36165),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__7181 (
            .O(N__36162),
            .I(N__36158));
    CascadeMux I__7180 (
            .O(N__36161),
            .I(N__36155));
    InMux I__7179 (
            .O(N__36158),
            .I(N__36150));
    InMux I__7178 (
            .O(N__36155),
            .I(N__36150));
    LocalMux I__7177 (
            .O(N__36150),
            .I(N__36146));
    InMux I__7176 (
            .O(N__36149),
            .I(N__36143));
    Span4Mux_h I__7175 (
            .O(N__36146),
            .I(N__36140));
    LocalMux I__7174 (
            .O(N__36143),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__7173 (
            .O(N__36140),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__7172 (
            .O(N__36135),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__7171 (
            .O(N__36132),
            .I(N__36128));
    CascadeMux I__7170 (
            .O(N__36131),
            .I(N__36125));
    InMux I__7169 (
            .O(N__36128),
            .I(N__36119));
    InMux I__7168 (
            .O(N__36125),
            .I(N__36119));
    InMux I__7167 (
            .O(N__36124),
            .I(N__36116));
    LocalMux I__7166 (
            .O(N__36119),
            .I(N__36113));
    LocalMux I__7165 (
            .O(N__36116),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__7164 (
            .O(N__36113),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__7163 (
            .O(N__36108),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__7162 (
            .O(N__36105),
            .I(N__36098));
    InMux I__7161 (
            .O(N__36104),
            .I(N__36098));
    InMux I__7160 (
            .O(N__36103),
            .I(N__36095));
    LocalMux I__7159 (
            .O(N__36098),
            .I(N__36092));
    LocalMux I__7158 (
            .O(N__36095),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__7157 (
            .O(N__36092),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__7156 (
            .O(N__36087),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    CascadeMux I__7155 (
            .O(N__36084),
            .I(N__36081));
    InMux I__7154 (
            .O(N__36081),
            .I(N__36077));
    InMux I__7153 (
            .O(N__36080),
            .I(N__36074));
    LocalMux I__7152 (
            .O(N__36077),
            .I(N__36068));
    LocalMux I__7151 (
            .O(N__36074),
            .I(N__36068));
    InMux I__7150 (
            .O(N__36073),
            .I(N__36065));
    Span4Mux_h I__7149 (
            .O(N__36068),
            .I(N__36062));
    LocalMux I__7148 (
            .O(N__36065),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__7147 (
            .O(N__36062),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__7146 (
            .O(N__36057),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__7145 (
            .O(N__36054),
            .I(N__36051));
    InMux I__7144 (
            .O(N__36051),
            .I(N__36046));
    CascadeMux I__7143 (
            .O(N__36050),
            .I(N__36043));
    InMux I__7142 (
            .O(N__36049),
            .I(N__36040));
    LocalMux I__7141 (
            .O(N__36046),
            .I(N__36037));
    InMux I__7140 (
            .O(N__36043),
            .I(N__36034));
    LocalMux I__7139 (
            .O(N__36040),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__7138 (
            .O(N__36037),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    LocalMux I__7137 (
            .O(N__36034),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__7136 (
            .O(N__36027),
            .I(bfn_14_7_0_));
    InMux I__7135 (
            .O(N__36024),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__7134 (
            .O(N__36021),
            .I(N__36017));
    CascadeMux I__7133 (
            .O(N__36020),
            .I(N__36014));
    InMux I__7132 (
            .O(N__36017),
            .I(N__36008));
    InMux I__7131 (
            .O(N__36014),
            .I(N__36008));
    InMux I__7130 (
            .O(N__36013),
            .I(N__36005));
    LocalMux I__7129 (
            .O(N__36008),
            .I(N__36002));
    LocalMux I__7128 (
            .O(N__36005),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv4 I__7127 (
            .O(N__36002),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__7126 (
            .O(N__35997),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    CascadeMux I__7125 (
            .O(N__35994),
            .I(N__35991));
    InMux I__7124 (
            .O(N__35991),
            .I(N__35987));
    InMux I__7123 (
            .O(N__35990),
            .I(N__35983));
    LocalMux I__7122 (
            .O(N__35987),
            .I(N__35980));
    InMux I__7121 (
            .O(N__35986),
            .I(N__35977));
    LocalMux I__7120 (
            .O(N__35983),
            .I(N__35974));
    Span4Mux_v I__7119 (
            .O(N__35980),
            .I(N__35971));
    LocalMux I__7118 (
            .O(N__35977),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__7117 (
            .O(N__35974),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__7116 (
            .O(N__35971),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__7115 (
            .O(N__35964),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__7114 (
            .O(N__35961),
            .I(N__35954));
    InMux I__7113 (
            .O(N__35960),
            .I(N__35954));
    InMux I__7112 (
            .O(N__35959),
            .I(N__35951));
    LocalMux I__7111 (
            .O(N__35954),
            .I(N__35948));
    LocalMux I__7110 (
            .O(N__35951),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__7109 (
            .O(N__35948),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__7108 (
            .O(N__35943),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__7107 (
            .O(N__35940),
            .I(N__35936));
    CascadeMux I__7106 (
            .O(N__35939),
            .I(N__35933));
    InMux I__7105 (
            .O(N__35936),
            .I(N__35927));
    InMux I__7104 (
            .O(N__35933),
            .I(N__35927));
    InMux I__7103 (
            .O(N__35932),
            .I(N__35924));
    LocalMux I__7102 (
            .O(N__35927),
            .I(N__35921));
    LocalMux I__7101 (
            .O(N__35924),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__7100 (
            .O(N__35921),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__7099 (
            .O(N__35916),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CascadeMux I__7098 (
            .O(N__35913),
            .I(N__35909));
    CascadeMux I__7097 (
            .O(N__35912),
            .I(N__35906));
    InMux I__7096 (
            .O(N__35909),
            .I(N__35901));
    InMux I__7095 (
            .O(N__35906),
            .I(N__35901));
    LocalMux I__7094 (
            .O(N__35901),
            .I(N__35897));
    InMux I__7093 (
            .O(N__35900),
            .I(N__35894));
    Span4Mux_h I__7092 (
            .O(N__35897),
            .I(N__35891));
    LocalMux I__7091 (
            .O(N__35894),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__7090 (
            .O(N__35891),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__7089 (
            .O(N__35886),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    CascadeMux I__7088 (
            .O(N__35883),
            .I(N__35879));
    InMux I__7087 (
            .O(N__35882),
            .I(N__35876));
    InMux I__7086 (
            .O(N__35879),
            .I(N__35872));
    LocalMux I__7085 (
            .O(N__35876),
            .I(N__35869));
    InMux I__7084 (
            .O(N__35875),
            .I(N__35866));
    LocalMux I__7083 (
            .O(N__35872),
            .I(N__35861));
    Span4Mux_h I__7082 (
            .O(N__35869),
            .I(N__35861));
    LocalMux I__7081 (
            .O(N__35866),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__7080 (
            .O(N__35861),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__7079 (
            .O(N__35856),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__7078 (
            .O(N__35853),
            .I(N__35850));
    InMux I__7077 (
            .O(N__35850),
            .I(N__35846));
    InMux I__7076 (
            .O(N__35849),
            .I(N__35842));
    LocalMux I__7075 (
            .O(N__35846),
            .I(N__35839));
    InMux I__7074 (
            .O(N__35845),
            .I(N__35836));
    LocalMux I__7073 (
            .O(N__35842),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__7072 (
            .O(N__35839),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    LocalMux I__7071 (
            .O(N__35836),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__7070 (
            .O(N__35829),
            .I(bfn_14_6_0_));
    IoInMux I__7069 (
            .O(N__35826),
            .I(N__35823));
    LocalMux I__7068 (
            .O(N__35823),
            .I(N__35820));
    Span12Mux_s1_v I__7067 (
            .O(N__35820),
            .I(N__35817));
    Odrv12 I__7066 (
            .O(N__35817),
            .I(\current_shift_inst.timer_s1.N_166_i ));
    InMux I__7065 (
            .O(N__35814),
            .I(N__35810));
    InMux I__7064 (
            .O(N__35813),
            .I(N__35807));
    LocalMux I__7063 (
            .O(N__35810),
            .I(N__35801));
    LocalMux I__7062 (
            .O(N__35807),
            .I(N__35801));
    InMux I__7061 (
            .O(N__35806),
            .I(N__35797));
    Span12Mux_s10_v I__7060 (
            .O(N__35801),
            .I(N__35794));
    InMux I__7059 (
            .O(N__35800),
            .I(N__35791));
    LocalMux I__7058 (
            .O(N__35797),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__7057 (
            .O(N__35794),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__7056 (
            .O(N__35791),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__7055 (
            .O(N__35784),
            .I(N__35781));
    LocalMux I__7054 (
            .O(N__35781),
            .I(N__35776));
    InMux I__7053 (
            .O(N__35780),
            .I(N__35770));
    InMux I__7052 (
            .O(N__35779),
            .I(N__35770));
    Span12Mux_s11_v I__7051 (
            .O(N__35776),
            .I(N__35767));
    InMux I__7050 (
            .O(N__35775),
            .I(N__35764));
    LocalMux I__7049 (
            .O(N__35770),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv12 I__7048 (
            .O(N__35767),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7047 (
            .O(N__35764),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    InMux I__7046 (
            .O(N__35757),
            .I(N__35754));
    LocalMux I__7045 (
            .O(N__35754),
            .I(N__35751));
    Span12Mux_s9_v I__7044 (
            .O(N__35751),
            .I(N__35745));
    InMux I__7043 (
            .O(N__35750),
            .I(N__35740));
    InMux I__7042 (
            .O(N__35749),
            .I(N__35740));
    InMux I__7041 (
            .O(N__35748),
            .I(N__35737));
    Span12Mux_v I__7040 (
            .O(N__35745),
            .I(N__35734));
    LocalMux I__7039 (
            .O(N__35740),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__7038 (
            .O(N__35737),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv12 I__7037 (
            .O(N__35734),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    IoInMux I__7036 (
            .O(N__35727),
            .I(N__35724));
    LocalMux I__7035 (
            .O(N__35724),
            .I(N__35720));
    InMux I__7034 (
            .O(N__35723),
            .I(N__35717));
    Span12Mux_s5_v I__7033 (
            .O(N__35720),
            .I(N__35713));
    LocalMux I__7032 (
            .O(N__35717),
            .I(N__35710));
    InMux I__7031 (
            .O(N__35716),
            .I(N__35707));
    Odrv12 I__7030 (
            .O(N__35713),
            .I(s1_phy_c));
    Odrv4 I__7029 (
            .O(N__35710),
            .I(s1_phy_c));
    LocalMux I__7028 (
            .O(N__35707),
            .I(s1_phy_c));
    IoInMux I__7027 (
            .O(N__35700),
            .I(N__35697));
    LocalMux I__7026 (
            .O(N__35697),
            .I(N__35694));
    Span4Mux_s2_v I__7025 (
            .O(N__35694),
            .I(N__35691));
    Span4Mux_h I__7024 (
            .O(N__35691),
            .I(N__35687));
    InMux I__7023 (
            .O(N__35690),
            .I(N__35684));
    Odrv4 I__7022 (
            .O(N__35687),
            .I(T23_c));
    LocalMux I__7021 (
            .O(N__35684),
            .I(T23_c));
    InMux I__7020 (
            .O(N__35679),
            .I(N__35673));
    InMux I__7019 (
            .O(N__35678),
            .I(N__35673));
    LocalMux I__7018 (
            .O(N__35673),
            .I(N__35670));
    Span4Mux_v I__7017 (
            .O(N__35670),
            .I(N__35665));
    InMux I__7016 (
            .O(N__35669),
            .I(N__35662));
    InMux I__7015 (
            .O(N__35668),
            .I(N__35659));
    Odrv4 I__7014 (
            .O(N__35665),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__7013 (
            .O(N__35662),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__7012 (
            .O(N__35659),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    CascadeMux I__7011 (
            .O(N__35652),
            .I(N__35646));
    InMux I__7010 (
            .O(N__35651),
            .I(N__35642));
    InMux I__7009 (
            .O(N__35650),
            .I(N__35639));
    InMux I__7008 (
            .O(N__35649),
            .I(N__35636));
    InMux I__7007 (
            .O(N__35646),
            .I(N__35633));
    InMux I__7006 (
            .O(N__35645),
            .I(N__35630));
    LocalMux I__7005 (
            .O(N__35642),
            .I(N__35625));
    LocalMux I__7004 (
            .O(N__35639),
            .I(N__35616));
    LocalMux I__7003 (
            .O(N__35636),
            .I(N__35616));
    LocalMux I__7002 (
            .O(N__35633),
            .I(N__35616));
    LocalMux I__7001 (
            .O(N__35630),
            .I(N__35616));
    InMux I__7000 (
            .O(N__35629),
            .I(N__35612));
    InMux I__6999 (
            .O(N__35628),
            .I(N__35609));
    Span4Mux_v I__6998 (
            .O(N__35625),
            .I(N__35604));
    Span4Mux_v I__6997 (
            .O(N__35616),
            .I(N__35604));
    InMux I__6996 (
            .O(N__35615),
            .I(N__35601));
    LocalMux I__6995 (
            .O(N__35612),
            .I(state_3));
    LocalMux I__6994 (
            .O(N__35609),
            .I(state_3));
    Odrv4 I__6993 (
            .O(N__35604),
            .I(state_3));
    LocalMux I__6992 (
            .O(N__35601),
            .I(state_3));
    IoInMux I__6991 (
            .O(N__35592),
            .I(N__35589));
    LocalMux I__6990 (
            .O(N__35589),
            .I(N__35586));
    Span4Mux_s0_v I__6989 (
            .O(N__35586),
            .I(N__35583));
    Span4Mux_v I__6988 (
            .O(N__35583),
            .I(N__35579));
    InMux I__6987 (
            .O(N__35582),
            .I(N__35576));
    Odrv4 I__6986 (
            .O(N__35579),
            .I(T45_c));
    LocalMux I__6985 (
            .O(N__35576),
            .I(T45_c));
    CascadeMux I__6984 (
            .O(N__35571),
            .I(N__35565));
    InMux I__6983 (
            .O(N__35570),
            .I(N__35561));
    InMux I__6982 (
            .O(N__35569),
            .I(N__35558));
    CascadeMux I__6981 (
            .O(N__35568),
            .I(N__35554));
    InMux I__6980 (
            .O(N__35565),
            .I(N__35551));
    InMux I__6979 (
            .O(N__35564),
            .I(N__35548));
    LocalMux I__6978 (
            .O(N__35561),
            .I(N__35545));
    LocalMux I__6977 (
            .O(N__35558),
            .I(N__35542));
    InMux I__6976 (
            .O(N__35557),
            .I(N__35539));
    InMux I__6975 (
            .O(N__35554),
            .I(N__35536));
    LocalMux I__6974 (
            .O(N__35551),
            .I(N__35533));
    LocalMux I__6973 (
            .O(N__35548),
            .I(N__35530));
    Span4Mux_h I__6972 (
            .O(N__35545),
            .I(N__35527));
    Span4Mux_h I__6971 (
            .O(N__35542),
            .I(N__35524));
    LocalMux I__6970 (
            .O(N__35539),
            .I(N__35521));
    LocalMux I__6969 (
            .O(N__35536),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__6968 (
            .O(N__35533),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__6967 (
            .O(N__35530),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__6966 (
            .O(N__35527),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__6965 (
            .O(N__35524),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__6964 (
            .O(N__35521),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__6963 (
            .O(N__35508),
            .I(N__35505));
    LocalMux I__6962 (
            .O(N__35505),
            .I(N__35502));
    Odrv12 I__6961 (
            .O(N__35502),
            .I(s2_phy_c));
    InMux I__6960 (
            .O(N__35499),
            .I(bfn_14_5_0_));
    CascadeMux I__6959 (
            .O(N__35496),
            .I(N__35493));
    InMux I__6958 (
            .O(N__35493),
            .I(N__35490));
    LocalMux I__6957 (
            .O(N__35490),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df22 ));
    InMux I__6956 (
            .O(N__35487),
            .I(N__35483));
    InMux I__6955 (
            .O(N__35486),
            .I(N__35480));
    LocalMux I__6954 (
            .O(N__35483),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    LocalMux I__6953 (
            .O(N__35480),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__6952 (
            .O(N__35475),
            .I(N__35471));
    InMux I__6951 (
            .O(N__35474),
            .I(N__35468));
    LocalMux I__6950 (
            .O(N__35471),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    LocalMux I__6949 (
            .O(N__35468),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__6948 (
            .O(N__35463),
            .I(N__35460));
    LocalMux I__6947 (
            .O(N__35460),
            .I(N__35457));
    Span4Mux_v I__6946 (
            .O(N__35457),
            .I(N__35454));
    Odrv4 I__6945 (
            .O(N__35454),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df20 ));
    InMux I__6944 (
            .O(N__35451),
            .I(N__35446));
    InMux I__6943 (
            .O(N__35450),
            .I(N__35443));
    InMux I__6942 (
            .O(N__35449),
            .I(N__35440));
    LocalMux I__6941 (
            .O(N__35446),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__6940 (
            .O(N__35443),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__6939 (
            .O(N__35440),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__6938 (
            .O(N__35433),
            .I(N__35430));
    LocalMux I__6937 (
            .O(N__35430),
            .I(N__35427));
    Odrv12 I__6936 (
            .O(N__35427),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    InMux I__6935 (
            .O(N__35424),
            .I(N__35420));
    InMux I__6934 (
            .O(N__35423),
            .I(N__35417));
    LocalMux I__6933 (
            .O(N__35420),
            .I(\phase_controller_inst1.time_passed_RNI7NN7 ));
    LocalMux I__6932 (
            .O(N__35417),
            .I(\phase_controller_inst1.time_passed_RNI7NN7 ));
    CascadeMux I__6931 (
            .O(N__35412),
            .I(N__35409));
    InMux I__6930 (
            .O(N__35409),
            .I(N__35404));
    InMux I__6929 (
            .O(N__35408),
            .I(N__35401));
    InMux I__6928 (
            .O(N__35407),
            .I(N__35397));
    LocalMux I__6927 (
            .O(N__35404),
            .I(N__35393));
    LocalMux I__6926 (
            .O(N__35401),
            .I(N__35390));
    InMux I__6925 (
            .O(N__35400),
            .I(N__35387));
    LocalMux I__6924 (
            .O(N__35397),
            .I(N__35384));
    InMux I__6923 (
            .O(N__35396),
            .I(N__35380));
    Span4Mux_h I__6922 (
            .O(N__35393),
            .I(N__35377));
    Span4Mux_h I__6921 (
            .O(N__35390),
            .I(N__35374));
    LocalMux I__6920 (
            .O(N__35387),
            .I(N__35369));
    Span12Mux_v I__6919 (
            .O(N__35384),
            .I(N__35369));
    InMux I__6918 (
            .O(N__35383),
            .I(N__35366));
    LocalMux I__6917 (
            .O(N__35380),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__6916 (
            .O(N__35377),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__6915 (
            .O(N__35374),
            .I(phase_controller_inst1_state_4));
    Odrv12 I__6914 (
            .O(N__35369),
            .I(phase_controller_inst1_state_4));
    LocalMux I__6913 (
            .O(N__35366),
            .I(phase_controller_inst1_state_4));
    InMux I__6912 (
            .O(N__35355),
            .I(N__35347));
    InMux I__6911 (
            .O(N__35354),
            .I(N__35347));
    InMux I__6910 (
            .O(N__35353),
            .I(N__35342));
    InMux I__6909 (
            .O(N__35352),
            .I(N__35342));
    LocalMux I__6908 (
            .O(N__35347),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__6907 (
            .O(N__35342),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__6906 (
            .O(N__35337),
            .I(N__35334));
    LocalMux I__6905 (
            .O(N__35334),
            .I(N__35331));
    Odrv12 I__6904 (
            .O(N__35331),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ));
    InMux I__6903 (
            .O(N__35328),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ));
    InMux I__6902 (
            .O(N__35325),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    InMux I__6901 (
            .O(N__35322),
            .I(N__35316));
    InMux I__6900 (
            .O(N__35321),
            .I(N__35316));
    LocalMux I__6899 (
            .O(N__35316),
            .I(N__35313));
    Odrv12 I__6898 (
            .O(N__35313),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__6897 (
            .O(N__35310),
            .I(N__35306));
    InMux I__6896 (
            .O(N__35309),
            .I(N__35303));
    LocalMux I__6895 (
            .O(N__35306),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    LocalMux I__6894 (
            .O(N__35303),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__6893 (
            .O(N__35298),
            .I(N__35294));
    InMux I__6892 (
            .O(N__35297),
            .I(N__35291));
    LocalMux I__6891 (
            .O(N__35294),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    LocalMux I__6890 (
            .O(N__35291),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__6889 (
            .O(N__35286),
            .I(N__35283));
    LocalMux I__6888 (
            .O(N__35283),
            .I(N__35280));
    Odrv4 I__6887 (
            .O(N__35280),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df22 ));
    InMux I__6886 (
            .O(N__35277),
            .I(N__35273));
    InMux I__6885 (
            .O(N__35276),
            .I(N__35270));
    LocalMux I__6884 (
            .O(N__35273),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__6883 (
            .O(N__35270),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__6882 (
            .O(N__35265),
            .I(N__35261));
    InMux I__6881 (
            .O(N__35264),
            .I(N__35258));
    LocalMux I__6880 (
            .O(N__35261),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__6879 (
            .O(N__35258),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    CascadeMux I__6878 (
            .O(N__35253),
            .I(N__35250));
    InMux I__6877 (
            .O(N__35250),
            .I(N__35247));
    LocalMux I__6876 (
            .O(N__35247),
            .I(N__35244));
    Odrv4 I__6875 (
            .O(N__35244),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df24 ));
    InMux I__6874 (
            .O(N__35241),
            .I(N__35237));
    InMux I__6873 (
            .O(N__35240),
            .I(N__35234));
    LocalMux I__6872 (
            .O(N__35237),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__6871 (
            .O(N__35234),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__6870 (
            .O(N__35229),
            .I(N__35225));
    InMux I__6869 (
            .O(N__35228),
            .I(N__35222));
    LocalMux I__6868 (
            .O(N__35225),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__6867 (
            .O(N__35222),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    CascadeMux I__6866 (
            .O(N__35217),
            .I(N__35214));
    InMux I__6865 (
            .O(N__35214),
            .I(N__35211));
    LocalMux I__6864 (
            .O(N__35211),
            .I(N__35208));
    Odrv4 I__6863 (
            .O(N__35208),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df26 ));
    InMux I__6862 (
            .O(N__35205),
            .I(N__35201));
    InMux I__6861 (
            .O(N__35204),
            .I(N__35198));
    LocalMux I__6860 (
            .O(N__35201),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__6859 (
            .O(N__35198),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__6858 (
            .O(N__35193),
            .I(N__35189));
    InMux I__6857 (
            .O(N__35192),
            .I(N__35186));
    LocalMux I__6856 (
            .O(N__35189),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__6855 (
            .O(N__35186),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__6854 (
            .O(N__35181),
            .I(N__35178));
    LocalMux I__6853 (
            .O(N__35178),
            .I(N__35175));
    Odrv4 I__6852 (
            .O(N__35175),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df28 ));
    InMux I__6851 (
            .O(N__35172),
            .I(N__35168));
    InMux I__6850 (
            .O(N__35171),
            .I(N__35165));
    LocalMux I__6849 (
            .O(N__35168),
            .I(N__35158));
    LocalMux I__6848 (
            .O(N__35165),
            .I(N__35158));
    InMux I__6847 (
            .O(N__35164),
            .I(N__35155));
    InMux I__6846 (
            .O(N__35163),
            .I(N__35152));
    Span4Mux_v I__6845 (
            .O(N__35158),
            .I(N__35149));
    LocalMux I__6844 (
            .O(N__35155),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    LocalMux I__6843 (
            .O(N__35152),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__6842 (
            .O(N__35149),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__6841 (
            .O(N__35142),
            .I(N__35139));
    LocalMux I__6840 (
            .O(N__35139),
            .I(N__35134));
    InMux I__6839 (
            .O(N__35138),
            .I(N__35131));
    InMux I__6838 (
            .O(N__35137),
            .I(N__35128));
    Span4Mux_h I__6837 (
            .O(N__35134),
            .I(N__35125));
    LocalMux I__6836 (
            .O(N__35131),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__6835 (
            .O(N__35128),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__6834 (
            .O(N__35125),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    CascadeMux I__6833 (
            .O(N__35118),
            .I(N__35115));
    InMux I__6832 (
            .O(N__35115),
            .I(N__35112));
    LocalMux I__6831 (
            .O(N__35112),
            .I(N__35109));
    Odrv4 I__6830 (
            .O(N__35109),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    InMux I__6829 (
            .O(N__35106),
            .I(N__35103));
    LocalMux I__6828 (
            .O(N__35103),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df20 ));
    CascadeMux I__6827 (
            .O(N__35100),
            .I(N__35097));
    InMux I__6826 (
            .O(N__35097),
            .I(N__35094));
    LocalMux I__6825 (
            .O(N__35094),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__6824 (
            .O(N__35091),
            .I(N__35088));
    LocalMux I__6823 (
            .O(N__35088),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__6822 (
            .O(N__35085),
            .I(N__35082));
    LocalMux I__6821 (
            .O(N__35082),
            .I(N__35079));
    Span4Mux_v I__6820 (
            .O(N__35079),
            .I(N__35076));
    Odrv4 I__6819 (
            .O(N__35076),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df26 ));
    InMux I__6818 (
            .O(N__35073),
            .I(N__35070));
    LocalMux I__6817 (
            .O(N__35070),
            .I(N__35067));
    Span4Mux_v I__6816 (
            .O(N__35067),
            .I(N__35064));
    Odrv4 I__6815 (
            .O(N__35064),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df28 ));
    InMux I__6814 (
            .O(N__35061),
            .I(N__35058));
    LocalMux I__6813 (
            .O(N__35058),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__6812 (
            .O(N__35055),
            .I(N__35052));
    InMux I__6811 (
            .O(N__35052),
            .I(N__35049));
    LocalMux I__6810 (
            .O(N__35049),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__6809 (
            .O(N__35046),
            .I(N__35043));
    InMux I__6808 (
            .O(N__35043),
            .I(N__35040));
    LocalMux I__6807 (
            .O(N__35040),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    CascadeMux I__6806 (
            .O(N__35037),
            .I(N__35034));
    InMux I__6805 (
            .O(N__35034),
            .I(N__35031));
    LocalMux I__6804 (
            .O(N__35031),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__6803 (
            .O(N__35028),
            .I(N__35025));
    InMux I__6802 (
            .O(N__35025),
            .I(N__35022));
    LocalMux I__6801 (
            .O(N__35022),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__6800 (
            .O(N__35019),
            .I(N__35016));
    InMux I__6799 (
            .O(N__35016),
            .I(N__35013));
    LocalMux I__6798 (
            .O(N__35013),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    CascadeMux I__6797 (
            .O(N__35010),
            .I(N__35007));
    InMux I__6796 (
            .O(N__35007),
            .I(N__35004));
    LocalMux I__6795 (
            .O(N__35004),
            .I(N__35001));
    Odrv4 I__6794 (
            .O(N__35001),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__6793 (
            .O(N__34998),
            .I(N__34995));
    InMux I__6792 (
            .O(N__34995),
            .I(N__34992));
    LocalMux I__6791 (
            .O(N__34992),
            .I(N__34989));
    Odrv4 I__6790 (
            .O(N__34989),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__6789 (
            .O(N__34986),
            .I(N__34981));
    InMux I__6788 (
            .O(N__34985),
            .I(N__34978));
    InMux I__6787 (
            .O(N__34984),
            .I(N__34975));
    LocalMux I__6786 (
            .O(N__34981),
            .I(N__34970));
    LocalMux I__6785 (
            .O(N__34978),
            .I(N__34970));
    LocalMux I__6784 (
            .O(N__34975),
            .I(\phase_controller_inst2.tr_time_passed ));
    Odrv12 I__6783 (
            .O(N__34970),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__6782 (
            .O(N__34965),
            .I(N__34959));
    InMux I__6781 (
            .O(N__34964),
            .I(N__34959));
    LocalMux I__6780 (
            .O(N__34959),
            .I(N__34954));
    CascadeMux I__6779 (
            .O(N__34958),
            .I(N__34951));
    InMux I__6778 (
            .O(N__34957),
            .I(N__34948));
    Span4Mux_h I__6777 (
            .O(N__34954),
            .I(N__34945));
    InMux I__6776 (
            .O(N__34951),
            .I(N__34942));
    LocalMux I__6775 (
            .O(N__34948),
            .I(N__34939));
    Span4Mux_h I__6774 (
            .O(N__34945),
            .I(N__34936));
    LocalMux I__6773 (
            .O(N__34942),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__6772 (
            .O(N__34939),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__6771 (
            .O(N__34936),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__6770 (
            .O(N__34929),
            .I(N__34926));
    LocalMux I__6769 (
            .O(N__34926),
            .I(N__34923));
    Span4Mux_h I__6768 (
            .O(N__34923),
            .I(N__34920));
    Span4Mux_h I__6767 (
            .O(N__34920),
            .I(N__34913));
    InMux I__6766 (
            .O(N__34919),
            .I(N__34904));
    InMux I__6765 (
            .O(N__34918),
            .I(N__34904));
    InMux I__6764 (
            .O(N__34917),
            .I(N__34904));
    InMux I__6763 (
            .O(N__34916),
            .I(N__34904));
    Odrv4 I__6762 (
            .O(N__34913),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__6761 (
            .O(N__34904),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    CascadeMux I__6760 (
            .O(N__34899),
            .I(N__34895));
    CascadeMux I__6759 (
            .O(N__34898),
            .I(N__34892));
    InMux I__6758 (
            .O(N__34895),
            .I(N__34884));
    InMux I__6757 (
            .O(N__34892),
            .I(N__34884));
    InMux I__6756 (
            .O(N__34891),
            .I(N__34881));
    InMux I__6755 (
            .O(N__34890),
            .I(N__34876));
    InMux I__6754 (
            .O(N__34889),
            .I(N__34876));
    LocalMux I__6753 (
            .O(N__34884),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__6752 (
            .O(N__34881),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__6751 (
            .O(N__34876),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__6750 (
            .O(N__34869),
            .I(N__34865));
    InMux I__6749 (
            .O(N__34868),
            .I(N__34862));
    LocalMux I__6748 (
            .O(N__34865),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__6747 (
            .O(N__34862),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__6746 (
            .O(N__34857),
            .I(N__34854));
    InMux I__6745 (
            .O(N__34854),
            .I(N__34851));
    LocalMux I__6744 (
            .O(N__34851),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__6743 (
            .O(N__34848),
            .I(N__34845));
    InMux I__6742 (
            .O(N__34845),
            .I(N__34842));
    LocalMux I__6741 (
            .O(N__34842),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    CascadeMux I__6740 (
            .O(N__34839),
            .I(N__34836));
    InMux I__6739 (
            .O(N__34836),
            .I(N__34833));
    LocalMux I__6738 (
            .O(N__34833),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__6737 (
            .O(N__34830),
            .I(N__34827));
    InMux I__6736 (
            .O(N__34827),
            .I(N__34824));
    LocalMux I__6735 (
            .O(N__34824),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    CascadeMux I__6734 (
            .O(N__34821),
            .I(N__34818));
    InMux I__6733 (
            .O(N__34818),
            .I(N__34815));
    LocalMux I__6732 (
            .O(N__34815),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__6731 (
            .O(N__34812),
            .I(N__34809));
    LocalMux I__6730 (
            .O(N__34809),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__6729 (
            .O(N__34806),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__6728 (
            .O(N__34803),
            .I(N__34800));
    LocalMux I__6727 (
            .O(N__34800),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__6726 (
            .O(N__34797),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__6725 (
            .O(N__34794),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__6724 (
            .O(N__34791),
            .I(N__34787));
    InMux I__6723 (
            .O(N__34790),
            .I(N__34784));
    LocalMux I__6722 (
            .O(N__34787),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__6721 (
            .O(N__34784),
            .I(\current_shift_inst.control_input_31 ));
    CascadeMux I__6720 (
            .O(N__34779),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__6719 (
            .O(N__34776),
            .I(N__34770));
    InMux I__6718 (
            .O(N__34775),
            .I(N__34770));
    LocalMux I__6717 (
            .O(N__34770),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__6716 (
            .O(N__34767),
            .I(N__34764));
    LocalMux I__6715 (
            .O(N__34764),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__6714 (
            .O(N__34761),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__6713 (
            .O(N__34758),
            .I(N__34755));
    LocalMux I__6712 (
            .O(N__34755),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__6711 (
            .O(N__34752),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__6710 (
            .O(N__34749),
            .I(N__34746));
    LocalMux I__6709 (
            .O(N__34746),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__6708 (
            .O(N__34743),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__6707 (
            .O(N__34740),
            .I(N__34737));
    LocalMux I__6706 (
            .O(N__34737),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__6705 (
            .O(N__34734),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__6704 (
            .O(N__34731),
            .I(N__34728));
    LocalMux I__6703 (
            .O(N__34728),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__6702 (
            .O(N__34725),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__6701 (
            .O(N__34722),
            .I(N__34719));
    LocalMux I__6700 (
            .O(N__34719),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__6699 (
            .O(N__34716),
            .I(bfn_13_12_0_));
    InMux I__6698 (
            .O(N__34713),
            .I(N__34710));
    LocalMux I__6697 (
            .O(N__34710),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__6696 (
            .O(N__34707),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__6695 (
            .O(N__34704),
            .I(N__34701));
    LocalMux I__6694 (
            .O(N__34701),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__6693 (
            .O(N__34698),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__6692 (
            .O(N__34695),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__6691 (
            .O(N__34692),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__6690 (
            .O(N__34689),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__6689 (
            .O(N__34686),
            .I(N__34683));
    LocalMux I__6688 (
            .O(N__34683),
            .I(\current_shift_inst.control_input_18 ));
    InMux I__6687 (
            .O(N__34680),
            .I(N__34677));
    LocalMux I__6686 (
            .O(N__34677),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__6685 (
            .O(N__34674),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__6684 (
            .O(N__34671),
            .I(N__34668));
    LocalMux I__6683 (
            .O(N__34668),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__6682 (
            .O(N__34665),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__6681 (
            .O(N__34662),
            .I(bfn_13_9_0_));
    InMux I__6680 (
            .O(N__34659),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__6679 (
            .O(N__34656),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__6678 (
            .O(N__34653),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__6677 (
            .O(N__34650),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__6676 (
            .O(N__34647),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__6675 (
            .O(N__34644),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__6674 (
            .O(N__34641),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__6673 (
            .O(N__34638),
            .I(bfn_13_10_0_));
    InMux I__6672 (
            .O(N__34635),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__6671 (
            .O(N__34632),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__6670 (
            .O(N__34629),
            .I(bfn_13_8_0_));
    InMux I__6669 (
            .O(N__34626),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__6668 (
            .O(N__34623),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__6667 (
            .O(N__34620),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__6666 (
            .O(N__34617),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__6665 (
            .O(N__34614),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__6664 (
            .O(N__34611),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__6663 (
            .O(N__34608),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__6662 (
            .O(N__34605),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__6661 (
            .O(N__34602),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__6660 (
            .O(N__34599),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__6659 (
            .O(N__34596),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__6658 (
            .O(N__34593),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__6657 (
            .O(N__34590),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__6656 (
            .O(N__34587),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__6655 (
            .O(N__34584),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__6654 (
            .O(N__34581),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__6653 (
            .O(N__34578),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    CEMux I__6652 (
            .O(N__34575),
            .I(N__34564));
    CEMux I__6651 (
            .O(N__34574),
            .I(N__34548));
    InMux I__6650 (
            .O(N__34573),
            .I(N__34541));
    InMux I__6649 (
            .O(N__34572),
            .I(N__34541));
    InMux I__6648 (
            .O(N__34571),
            .I(N__34541));
    InMux I__6647 (
            .O(N__34570),
            .I(N__34532));
    InMux I__6646 (
            .O(N__34569),
            .I(N__34532));
    InMux I__6645 (
            .O(N__34568),
            .I(N__34532));
    InMux I__6644 (
            .O(N__34567),
            .I(N__34532));
    LocalMux I__6643 (
            .O(N__34564),
            .I(N__34525));
    InMux I__6642 (
            .O(N__34563),
            .I(N__34516));
    InMux I__6641 (
            .O(N__34562),
            .I(N__34516));
    InMux I__6640 (
            .O(N__34561),
            .I(N__34516));
    InMux I__6639 (
            .O(N__34560),
            .I(N__34516));
    CEMux I__6638 (
            .O(N__34559),
            .I(N__34503));
    CEMux I__6637 (
            .O(N__34558),
            .I(N__34499));
    InMux I__6636 (
            .O(N__34557),
            .I(N__34492));
    InMux I__6635 (
            .O(N__34556),
            .I(N__34492));
    InMux I__6634 (
            .O(N__34555),
            .I(N__34492));
    InMux I__6633 (
            .O(N__34554),
            .I(N__34483));
    InMux I__6632 (
            .O(N__34553),
            .I(N__34483));
    InMux I__6631 (
            .O(N__34552),
            .I(N__34483));
    InMux I__6630 (
            .O(N__34551),
            .I(N__34483));
    LocalMux I__6629 (
            .O(N__34548),
            .I(N__34480));
    LocalMux I__6628 (
            .O(N__34541),
            .I(N__34477));
    LocalMux I__6627 (
            .O(N__34532),
            .I(N__34474));
    InMux I__6626 (
            .O(N__34531),
            .I(N__34465));
    InMux I__6625 (
            .O(N__34530),
            .I(N__34465));
    InMux I__6624 (
            .O(N__34529),
            .I(N__34465));
    InMux I__6623 (
            .O(N__34528),
            .I(N__34465));
    Span4Mux_h I__6622 (
            .O(N__34525),
            .I(N__34460));
    LocalMux I__6621 (
            .O(N__34516),
            .I(N__34460));
    InMux I__6620 (
            .O(N__34515),
            .I(N__34451));
    InMux I__6619 (
            .O(N__34514),
            .I(N__34451));
    InMux I__6618 (
            .O(N__34513),
            .I(N__34451));
    InMux I__6617 (
            .O(N__34512),
            .I(N__34451));
    InMux I__6616 (
            .O(N__34511),
            .I(N__34442));
    InMux I__6615 (
            .O(N__34510),
            .I(N__34442));
    InMux I__6614 (
            .O(N__34509),
            .I(N__34442));
    InMux I__6613 (
            .O(N__34508),
            .I(N__34442));
    CEMux I__6612 (
            .O(N__34507),
            .I(N__34438));
    CEMux I__6611 (
            .O(N__34506),
            .I(N__34435));
    LocalMux I__6610 (
            .O(N__34503),
            .I(N__34432));
    CEMux I__6609 (
            .O(N__34502),
            .I(N__34429));
    LocalMux I__6608 (
            .O(N__34499),
            .I(N__34426));
    LocalMux I__6607 (
            .O(N__34492),
            .I(N__34407));
    LocalMux I__6606 (
            .O(N__34483),
            .I(N__34407));
    Span4Mux_v I__6605 (
            .O(N__34480),
            .I(N__34407));
    Span4Mux_v I__6604 (
            .O(N__34477),
            .I(N__34407));
    Span4Mux_h I__6603 (
            .O(N__34474),
            .I(N__34407));
    LocalMux I__6602 (
            .O(N__34465),
            .I(N__34407));
    Span4Mux_v I__6601 (
            .O(N__34460),
            .I(N__34407));
    LocalMux I__6600 (
            .O(N__34451),
            .I(N__34407));
    LocalMux I__6599 (
            .O(N__34442),
            .I(N__34407));
    InMux I__6598 (
            .O(N__34441),
            .I(N__34404));
    LocalMux I__6597 (
            .O(N__34438),
            .I(N__34401));
    LocalMux I__6596 (
            .O(N__34435),
            .I(N__34396));
    Span4Mux_h I__6595 (
            .O(N__34432),
            .I(N__34396));
    LocalMux I__6594 (
            .O(N__34429),
            .I(N__34391));
    Span4Mux_h I__6593 (
            .O(N__34426),
            .I(N__34391));
    Span4Mux_v I__6592 (
            .O(N__34407),
            .I(N__34386));
    LocalMux I__6591 (
            .O(N__34404),
            .I(N__34386));
    Span4Mux_h I__6590 (
            .O(N__34401),
            .I(N__34383));
    Span4Mux_h I__6589 (
            .O(N__34396),
            .I(N__34378));
    Span4Mux_h I__6588 (
            .O(N__34391),
            .I(N__34378));
    Span4Mux_h I__6587 (
            .O(N__34386),
            .I(N__34375));
    Odrv4 I__6586 (
            .O(N__34383),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__6585 (
            .O(N__34378),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__6584 (
            .O(N__34375),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__6583 (
            .O(N__34368),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__6582 (
            .O(N__34365),
            .I(N__34362));
    LocalMux I__6581 (
            .O(N__34362),
            .I(N__34358));
    InMux I__6580 (
            .O(N__34361),
            .I(N__34354));
    Span4Mux_h I__6579 (
            .O(N__34358),
            .I(N__34351));
    InMux I__6578 (
            .O(N__34357),
            .I(N__34348));
    LocalMux I__6577 (
            .O(N__34354),
            .I(N__34341));
    Sp12to4 I__6576 (
            .O(N__34351),
            .I(N__34341));
    LocalMux I__6575 (
            .O(N__34348),
            .I(N__34341));
    Span12Mux_s10_v I__6574 (
            .O(N__34341),
            .I(N__34338));
    Odrv12 I__6573 (
            .O(N__34338),
            .I(il_min_comp1_D2));
    IoInMux I__6572 (
            .O(N__34335),
            .I(N__34332));
    LocalMux I__6571 (
            .O(N__34332),
            .I(N__34329));
    IoSpan4Mux I__6570 (
            .O(N__34329),
            .I(N__34326));
    Span4Mux_s0_v I__6569 (
            .O(N__34326),
            .I(N__34323));
    Span4Mux_v I__6568 (
            .O(N__34323),
            .I(N__34319));
    InMux I__6567 (
            .O(N__34322),
            .I(N__34316));
    Odrv4 I__6566 (
            .O(N__34319),
            .I(T12_c));
    LocalMux I__6565 (
            .O(N__34316),
            .I(T12_c));
    InMux I__6564 (
            .O(N__34311),
            .I(N__34303));
    InMux I__6563 (
            .O(N__34310),
            .I(N__34303));
    InMux I__6562 (
            .O(N__34309),
            .I(N__34299));
    InMux I__6561 (
            .O(N__34308),
            .I(N__34296));
    LocalMux I__6560 (
            .O(N__34303),
            .I(N__34293));
    InMux I__6559 (
            .O(N__34302),
            .I(N__34290));
    LocalMux I__6558 (
            .O(N__34299),
            .I(N__34287));
    LocalMux I__6557 (
            .O(N__34296),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__6556 (
            .O(N__34293),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__6555 (
            .O(N__34290),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__6554 (
            .O(N__34287),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    IoInMux I__6553 (
            .O(N__34278),
            .I(N__34275));
    LocalMux I__6552 (
            .O(N__34275),
            .I(N__34272));
    Span4Mux_s0_v I__6551 (
            .O(N__34272),
            .I(N__34269));
    Span4Mux_v I__6550 (
            .O(N__34269),
            .I(N__34266));
    Sp12to4 I__6549 (
            .O(N__34266),
            .I(N__34262));
    InMux I__6548 (
            .O(N__34265),
            .I(N__34259));
    Odrv12 I__6547 (
            .O(N__34262),
            .I(T01_c));
    LocalMux I__6546 (
            .O(N__34259),
            .I(T01_c));
    CascadeMux I__6545 (
            .O(N__34254),
            .I(N__34250));
    InMux I__6544 (
            .O(N__34253),
            .I(N__34247));
    InMux I__6543 (
            .O(N__34250),
            .I(N__34243));
    LocalMux I__6542 (
            .O(N__34247),
            .I(N__34240));
    InMux I__6541 (
            .O(N__34246),
            .I(N__34237));
    LocalMux I__6540 (
            .O(N__34243),
            .I(N__34232));
    Span4Mux_h I__6539 (
            .O(N__34240),
            .I(N__34232));
    LocalMux I__6538 (
            .O(N__34237),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__6537 (
            .O(N__34232),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__6536 (
            .O(N__34227),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    CascadeMux I__6535 (
            .O(N__34224),
            .I(N__34221));
    InMux I__6534 (
            .O(N__34221),
            .I(N__34218));
    LocalMux I__6533 (
            .O(N__34218),
            .I(N__34213));
    InMux I__6532 (
            .O(N__34217),
            .I(N__34210));
    InMux I__6531 (
            .O(N__34216),
            .I(N__34207));
    Span4Mux_v I__6530 (
            .O(N__34213),
            .I(N__34204));
    LocalMux I__6529 (
            .O(N__34210),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__6528 (
            .O(N__34207),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__6527 (
            .O(N__34204),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__6526 (
            .O(N__34197),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__6525 (
            .O(N__34194),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__6524 (
            .O(N__34191),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__6523 (
            .O(N__34188),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__6522 (
            .O(N__34185),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__6521 (
            .O(N__34182),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__6520 (
            .O(N__34179),
            .I(bfn_12_20_0_));
    InMux I__6519 (
            .O(N__34176),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__6518 (
            .O(N__34173),
            .I(N__34169));
    InMux I__6517 (
            .O(N__34172),
            .I(N__34166));
    LocalMux I__6516 (
            .O(N__34169),
            .I(N__34163));
    LocalMux I__6515 (
            .O(N__34166),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__6514 (
            .O(N__34163),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__6513 (
            .O(N__34158),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__6512 (
            .O(N__34155),
            .I(N__34151));
    InMux I__6511 (
            .O(N__34154),
            .I(N__34148));
    LocalMux I__6510 (
            .O(N__34151),
            .I(N__34145));
    LocalMux I__6509 (
            .O(N__34148),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__6508 (
            .O(N__34145),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__6507 (
            .O(N__34140),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__6506 (
            .O(N__34137),
            .I(N__34133));
    InMux I__6505 (
            .O(N__34136),
            .I(N__34130));
    LocalMux I__6504 (
            .O(N__34133),
            .I(N__34127));
    LocalMux I__6503 (
            .O(N__34130),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__6502 (
            .O(N__34127),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__6501 (
            .O(N__34122),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__6500 (
            .O(N__34119),
            .I(N__34115));
    InMux I__6499 (
            .O(N__34118),
            .I(N__34112));
    LocalMux I__6498 (
            .O(N__34115),
            .I(N__34109));
    LocalMux I__6497 (
            .O(N__34112),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__6496 (
            .O(N__34109),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__6495 (
            .O(N__34104),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__6494 (
            .O(N__34101),
            .I(N__34097));
    InMux I__6493 (
            .O(N__34100),
            .I(N__34094));
    LocalMux I__6492 (
            .O(N__34097),
            .I(N__34091));
    LocalMux I__6491 (
            .O(N__34094),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__6490 (
            .O(N__34091),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__6489 (
            .O(N__34086),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__6488 (
            .O(N__34083),
            .I(N__34079));
    InMux I__6487 (
            .O(N__34082),
            .I(N__34076));
    LocalMux I__6486 (
            .O(N__34079),
            .I(N__34073));
    LocalMux I__6485 (
            .O(N__34076),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv12 I__6484 (
            .O(N__34073),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__6483 (
            .O(N__34068),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    CascadeMux I__6482 (
            .O(N__34065),
            .I(N__34061));
    InMux I__6481 (
            .O(N__34064),
            .I(N__34056));
    InMux I__6480 (
            .O(N__34061),
            .I(N__34056));
    LocalMux I__6479 (
            .O(N__34056),
            .I(N__34052));
    InMux I__6478 (
            .O(N__34055),
            .I(N__34049));
    Span4Mux_h I__6477 (
            .O(N__34052),
            .I(N__34046));
    LocalMux I__6476 (
            .O(N__34049),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__6475 (
            .O(N__34046),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__6474 (
            .O(N__34041),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    CascadeMux I__6473 (
            .O(N__34038),
            .I(N__34034));
    InMux I__6472 (
            .O(N__34037),
            .I(N__34029));
    InMux I__6471 (
            .O(N__34034),
            .I(N__34029));
    LocalMux I__6470 (
            .O(N__34029),
            .I(N__34025));
    InMux I__6469 (
            .O(N__34028),
            .I(N__34022));
    Span4Mux_h I__6468 (
            .O(N__34025),
            .I(N__34019));
    LocalMux I__6467 (
            .O(N__34022),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__6466 (
            .O(N__34019),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__6465 (
            .O(N__34014),
            .I(bfn_12_19_0_));
    CascadeMux I__6464 (
            .O(N__34011),
            .I(N__34008));
    InMux I__6463 (
            .O(N__34008),
            .I(N__34005));
    LocalMux I__6462 (
            .O(N__34005),
            .I(N__34002));
    Odrv4 I__6461 (
            .O(N__34002),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    InMux I__6460 (
            .O(N__33999),
            .I(N__33995));
    InMux I__6459 (
            .O(N__33998),
            .I(N__33992));
    LocalMux I__6458 (
            .O(N__33995),
            .I(N__33989));
    LocalMux I__6457 (
            .O(N__33992),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__6456 (
            .O(N__33989),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__6455 (
            .O(N__33984),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__6454 (
            .O(N__33981),
            .I(N__33978));
    LocalMux I__6453 (
            .O(N__33978),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28 ));
    CascadeMux I__6452 (
            .O(N__33975),
            .I(N__33971));
    InMux I__6451 (
            .O(N__33974),
            .I(N__33968));
    InMux I__6450 (
            .O(N__33971),
            .I(N__33965));
    LocalMux I__6449 (
            .O(N__33968),
            .I(N__33962));
    LocalMux I__6448 (
            .O(N__33965),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__6447 (
            .O(N__33962),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__6446 (
            .O(N__33957),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__6445 (
            .O(N__33954),
            .I(N__33950));
    InMux I__6444 (
            .O(N__33953),
            .I(N__33947));
    LocalMux I__6443 (
            .O(N__33950),
            .I(N__33944));
    LocalMux I__6442 (
            .O(N__33947),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__6441 (
            .O(N__33944),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__6440 (
            .O(N__33939),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__6439 (
            .O(N__33936),
            .I(N__33932));
    InMux I__6438 (
            .O(N__33935),
            .I(N__33929));
    LocalMux I__6437 (
            .O(N__33932),
            .I(N__33926));
    LocalMux I__6436 (
            .O(N__33929),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__6435 (
            .O(N__33926),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__6434 (
            .O(N__33921),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__6433 (
            .O(N__33918),
            .I(N__33914));
    InMux I__6432 (
            .O(N__33917),
            .I(N__33911));
    LocalMux I__6431 (
            .O(N__33914),
            .I(N__33908));
    LocalMux I__6430 (
            .O(N__33911),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__6429 (
            .O(N__33908),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__6428 (
            .O(N__33903),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__6427 (
            .O(N__33900),
            .I(N__33896));
    InMux I__6426 (
            .O(N__33899),
            .I(N__33893));
    LocalMux I__6425 (
            .O(N__33896),
            .I(N__33890));
    LocalMux I__6424 (
            .O(N__33893),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv12 I__6423 (
            .O(N__33890),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__6422 (
            .O(N__33885),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__6421 (
            .O(N__33882),
            .I(N__33879));
    LocalMux I__6420 (
            .O(N__33879),
            .I(N__33875));
    InMux I__6419 (
            .O(N__33878),
            .I(N__33872));
    Span4Mux_v I__6418 (
            .O(N__33875),
            .I(N__33869));
    LocalMux I__6417 (
            .O(N__33872),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__6416 (
            .O(N__33869),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__6415 (
            .O(N__33864),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__6414 (
            .O(N__33861),
            .I(N__33858));
    LocalMux I__6413 (
            .O(N__33858),
            .I(N__33854));
    InMux I__6412 (
            .O(N__33857),
            .I(N__33851));
    Span4Mux_v I__6411 (
            .O(N__33854),
            .I(N__33848));
    LocalMux I__6410 (
            .O(N__33851),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__6409 (
            .O(N__33848),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__6408 (
            .O(N__33843),
            .I(bfn_12_18_0_));
    InMux I__6407 (
            .O(N__33840),
            .I(N__33837));
    LocalMux I__6406 (
            .O(N__33837),
            .I(N__33834));
    Odrv4 I__6405 (
            .O(N__33834),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    CascadeMux I__6404 (
            .O(N__33831),
            .I(N__33828));
    InMux I__6403 (
            .O(N__33828),
            .I(N__33825));
    LocalMux I__6402 (
            .O(N__33825),
            .I(N__33822));
    Odrv12 I__6401 (
            .O(N__33822),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    CascadeMux I__6400 (
            .O(N__33819),
            .I(N__33816));
    InMux I__6399 (
            .O(N__33816),
            .I(N__33813));
    LocalMux I__6398 (
            .O(N__33813),
            .I(N__33810));
    Odrv12 I__6397 (
            .O(N__33810),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__6396 (
            .O(N__33807),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ));
    InMux I__6395 (
            .O(N__33804),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    InMux I__6394 (
            .O(N__33801),
            .I(N__33795));
    InMux I__6393 (
            .O(N__33800),
            .I(N__33795));
    LocalMux I__6392 (
            .O(N__33795),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    CascadeMux I__6391 (
            .O(N__33792),
            .I(N__33788));
    InMux I__6390 (
            .O(N__33791),
            .I(N__33785));
    InMux I__6389 (
            .O(N__33788),
            .I(N__33781));
    LocalMux I__6388 (
            .O(N__33785),
            .I(N__33778));
    InMux I__6387 (
            .O(N__33784),
            .I(N__33775));
    LocalMux I__6386 (
            .O(N__33781),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__6385 (
            .O(N__33778),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__6384 (
            .O(N__33775),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__6383 (
            .O(N__33768),
            .I(N__33765));
    LocalMux I__6382 (
            .O(N__33765),
            .I(N__33762));
    Span4Mux_h I__6381 (
            .O(N__33762),
            .I(N__33759));
    Odrv4 I__6380 (
            .O(N__33759),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__6379 (
            .O(N__33756),
            .I(N__33753));
    InMux I__6378 (
            .O(N__33753),
            .I(N__33750));
    LocalMux I__6377 (
            .O(N__33750),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__6376 (
            .O(N__33747),
            .I(N__33744));
    LocalMux I__6375 (
            .O(N__33744),
            .I(N__33741));
    Odrv4 I__6374 (
            .O(N__33741),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__6373 (
            .O(N__33738),
            .I(N__33735));
    InMux I__6372 (
            .O(N__33735),
            .I(N__33732));
    LocalMux I__6371 (
            .O(N__33732),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__6370 (
            .O(N__33729),
            .I(N__33726));
    InMux I__6369 (
            .O(N__33726),
            .I(N__33723));
    LocalMux I__6368 (
            .O(N__33723),
            .I(N__33720));
    Odrv4 I__6367 (
            .O(N__33720),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    InMux I__6366 (
            .O(N__33717),
            .I(N__33714));
    LocalMux I__6365 (
            .O(N__33714),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__6364 (
            .O(N__33711),
            .I(N__33708));
    LocalMux I__6363 (
            .O(N__33708),
            .I(N__33705));
    Odrv4 I__6362 (
            .O(N__33705),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    CascadeMux I__6361 (
            .O(N__33702),
            .I(N__33699));
    InMux I__6360 (
            .O(N__33699),
            .I(N__33696));
    LocalMux I__6359 (
            .O(N__33696),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__6358 (
            .O(N__33693),
            .I(N__33690));
    InMux I__6357 (
            .O(N__33690),
            .I(N__33687));
    LocalMux I__6356 (
            .O(N__33687),
            .I(N__33684));
    Odrv4 I__6355 (
            .O(N__33684),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__6354 (
            .O(N__33681),
            .I(N__33678));
    LocalMux I__6353 (
            .O(N__33678),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__6352 (
            .O(N__33675),
            .I(N__33672));
    LocalMux I__6351 (
            .O(N__33672),
            .I(N__33669));
    Span4Mux_h I__6350 (
            .O(N__33669),
            .I(N__33666));
    Span4Mux_v I__6349 (
            .O(N__33666),
            .I(N__33663));
    Odrv4 I__6348 (
            .O(N__33663),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__6347 (
            .O(N__33660),
            .I(N__33657));
    InMux I__6346 (
            .O(N__33657),
            .I(N__33654));
    LocalMux I__6345 (
            .O(N__33654),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__6344 (
            .O(N__33651),
            .I(N__33648));
    LocalMux I__6343 (
            .O(N__33648),
            .I(N__33645));
    Span4Mux_h I__6342 (
            .O(N__33645),
            .I(N__33642));
    Odrv4 I__6341 (
            .O(N__33642),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__6340 (
            .O(N__33639),
            .I(N__33636));
    InMux I__6339 (
            .O(N__33636),
            .I(N__33633));
    LocalMux I__6338 (
            .O(N__33633),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__6337 (
            .O(N__33630),
            .I(N__33627));
    LocalMux I__6336 (
            .O(N__33627),
            .I(N__33624));
    Span4Mux_v I__6335 (
            .O(N__33624),
            .I(N__33621));
    Odrv4 I__6334 (
            .O(N__33621),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    CascadeMux I__6333 (
            .O(N__33618),
            .I(N__33615));
    InMux I__6332 (
            .O(N__33615),
            .I(N__33612));
    LocalMux I__6331 (
            .O(N__33612),
            .I(N__33609));
    Span4Mux_v I__6330 (
            .O(N__33609),
            .I(N__33606));
    Odrv4 I__6329 (
            .O(N__33606),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    InMux I__6328 (
            .O(N__33603),
            .I(N__33600));
    LocalMux I__6327 (
            .O(N__33600),
            .I(N__33597));
    Odrv4 I__6326 (
            .O(N__33597),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__6325 (
            .O(N__33594),
            .I(N__33591));
    InMux I__6324 (
            .O(N__33591),
            .I(N__33588));
    LocalMux I__6323 (
            .O(N__33588),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__6322 (
            .O(N__33585),
            .I(N__33582));
    LocalMux I__6321 (
            .O(N__33582),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__6320 (
            .O(N__33579),
            .I(N__33576));
    InMux I__6319 (
            .O(N__33576),
            .I(N__33573));
    LocalMux I__6318 (
            .O(N__33573),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    InMux I__6317 (
            .O(N__33570),
            .I(N__33567));
    LocalMux I__6316 (
            .O(N__33567),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__6315 (
            .O(N__33564),
            .I(N__33561));
    InMux I__6314 (
            .O(N__33561),
            .I(N__33558));
    LocalMux I__6313 (
            .O(N__33558),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__6312 (
            .O(N__33555),
            .I(N__33552));
    LocalMux I__6311 (
            .O(N__33552),
            .I(N__33549));
    Odrv4 I__6310 (
            .O(N__33549),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__6309 (
            .O(N__33546),
            .I(N__33543));
    InMux I__6308 (
            .O(N__33543),
            .I(N__33540));
    LocalMux I__6307 (
            .O(N__33540),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__6306 (
            .O(N__33537),
            .I(N__33534));
    LocalMux I__6305 (
            .O(N__33534),
            .I(N__33531));
    Span4Mux_h I__6304 (
            .O(N__33531),
            .I(N__33528));
    Span4Mux_h I__6303 (
            .O(N__33528),
            .I(N__33525));
    Odrv4 I__6302 (
            .O(N__33525),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__6301 (
            .O(N__33522),
            .I(N__33519));
    InMux I__6300 (
            .O(N__33519),
            .I(N__33516));
    LocalMux I__6299 (
            .O(N__33516),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__6298 (
            .O(N__33513),
            .I(N__33510));
    InMux I__6297 (
            .O(N__33510),
            .I(N__33507));
    LocalMux I__6296 (
            .O(N__33507),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    InMux I__6295 (
            .O(N__33504),
            .I(N__33501));
    LocalMux I__6294 (
            .O(N__33501),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__6293 (
            .O(N__33498),
            .I(N__33495));
    LocalMux I__6292 (
            .O(N__33495),
            .I(N__33492));
    Span4Mux_h I__6291 (
            .O(N__33492),
            .I(N__33489));
    Span4Mux_v I__6290 (
            .O(N__33489),
            .I(N__33486));
    Odrv4 I__6289 (
            .O(N__33486),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__6288 (
            .O(N__33483),
            .I(N__33480));
    InMux I__6287 (
            .O(N__33480),
            .I(N__33477));
    LocalMux I__6286 (
            .O(N__33477),
            .I(N__33474));
    Odrv4 I__6285 (
            .O(N__33474),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__6284 (
            .O(N__33471),
            .I(N__33468));
    LocalMux I__6283 (
            .O(N__33468),
            .I(N__33465));
    Span4Mux_v I__6282 (
            .O(N__33465),
            .I(N__33462));
    Odrv4 I__6281 (
            .O(N__33462),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__6280 (
            .O(N__33459),
            .I(N__33456));
    InMux I__6279 (
            .O(N__33456),
            .I(N__33453));
    LocalMux I__6278 (
            .O(N__33453),
            .I(N__33450));
    Odrv4 I__6277 (
            .O(N__33450),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__6276 (
            .O(N__33447),
            .I(N__33444));
    LocalMux I__6275 (
            .O(N__33444),
            .I(N__33440));
    InMux I__6274 (
            .O(N__33443),
            .I(N__33437));
    Span4Mux_v I__6273 (
            .O(N__33440),
            .I(N__33432));
    LocalMux I__6272 (
            .O(N__33437),
            .I(N__33432));
    Span4Mux_h I__6271 (
            .O(N__33432),
            .I(N__33428));
    InMux I__6270 (
            .O(N__33431),
            .I(N__33425));
    Odrv4 I__6269 (
            .O(N__33428),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    LocalMux I__6268 (
            .O(N__33425),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__6267 (
            .O(N__33420),
            .I(N__33417));
    LocalMux I__6266 (
            .O(N__33417),
            .I(N__33414));
    Span4Mux_v I__6265 (
            .O(N__33414),
            .I(N__33411));
    Odrv4 I__6264 (
            .O(N__33411),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ));
    InMux I__6263 (
            .O(N__33408),
            .I(N__33405));
    LocalMux I__6262 (
            .O(N__33405),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    CascadeMux I__6261 (
            .O(N__33402),
            .I(N__33399));
    InMux I__6260 (
            .O(N__33399),
            .I(N__33396));
    LocalMux I__6259 (
            .O(N__33396),
            .I(N__33393));
    Odrv4 I__6258 (
            .O(N__33393),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ));
    CascadeMux I__6257 (
            .O(N__33390),
            .I(N__33387));
    InMux I__6256 (
            .O(N__33387),
            .I(N__33384));
    LocalMux I__6255 (
            .O(N__33384),
            .I(N__33381));
    Span4Mux_h I__6254 (
            .O(N__33381),
            .I(N__33376));
    InMux I__6253 (
            .O(N__33380),
            .I(N__33371));
    InMux I__6252 (
            .O(N__33379),
            .I(N__33371));
    Odrv4 I__6251 (
            .O(N__33376),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    LocalMux I__6250 (
            .O(N__33371),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__6249 (
            .O(N__33366),
            .I(N__33363));
    LocalMux I__6248 (
            .O(N__33363),
            .I(N__33360));
    Span4Mux_h I__6247 (
            .O(N__33360),
            .I(N__33357));
    Span4Mux_h I__6246 (
            .O(N__33357),
            .I(N__33354));
    Odrv4 I__6245 (
            .O(N__33354),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__6244 (
            .O(N__33351),
            .I(N__33348));
    LocalMux I__6243 (
            .O(N__33348),
            .I(N__33344));
    InMux I__6242 (
            .O(N__33347),
            .I(N__33341));
    Span12Mux_s10_v I__6241 (
            .O(N__33344),
            .I(N__33335));
    LocalMux I__6240 (
            .O(N__33341),
            .I(N__33335));
    InMux I__6239 (
            .O(N__33340),
            .I(N__33332));
    Odrv12 I__6238 (
            .O(N__33335),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    LocalMux I__6237 (
            .O(N__33332),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__6236 (
            .O(N__33327),
            .I(N__33324));
    LocalMux I__6235 (
            .O(N__33324),
            .I(N__33321));
    Span4Mux_h I__6234 (
            .O(N__33321),
            .I(N__33318));
    Odrv4 I__6233 (
            .O(N__33318),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ));
    CascadeMux I__6232 (
            .O(N__33315),
            .I(N__33311));
    InMux I__6231 (
            .O(N__33314),
            .I(N__33301));
    InMux I__6230 (
            .O(N__33311),
            .I(N__33301));
    InMux I__6229 (
            .O(N__33310),
            .I(N__33298));
    CascadeMux I__6228 (
            .O(N__33309),
            .I(N__33295));
    InMux I__6227 (
            .O(N__33308),
            .I(N__33288));
    InMux I__6226 (
            .O(N__33307),
            .I(N__33283));
    InMux I__6225 (
            .O(N__33306),
            .I(N__33283));
    LocalMux I__6224 (
            .O(N__33301),
            .I(N__33278));
    LocalMux I__6223 (
            .O(N__33298),
            .I(N__33278));
    InMux I__6222 (
            .O(N__33295),
            .I(N__33275));
    InMux I__6221 (
            .O(N__33294),
            .I(N__33270));
    InMux I__6220 (
            .O(N__33293),
            .I(N__33270));
    InMux I__6219 (
            .O(N__33292),
            .I(N__33267));
    InMux I__6218 (
            .O(N__33291),
            .I(N__33264));
    LocalMux I__6217 (
            .O(N__33288),
            .I(N__33257));
    LocalMux I__6216 (
            .O(N__33283),
            .I(N__33257));
    Span4Mux_v I__6215 (
            .O(N__33278),
            .I(N__33257));
    LocalMux I__6214 (
            .O(N__33275),
            .I(N__33252));
    LocalMux I__6213 (
            .O(N__33270),
            .I(N__33252));
    LocalMux I__6212 (
            .O(N__33267),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    LocalMux I__6211 (
            .O(N__33264),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    Odrv4 I__6210 (
            .O(N__33257),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    Odrv4 I__6209 (
            .O(N__33252),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    InMux I__6208 (
            .O(N__33243),
            .I(N__33231));
    InMux I__6207 (
            .O(N__33242),
            .I(N__33216));
    InMux I__6206 (
            .O(N__33241),
            .I(N__33216));
    InMux I__6205 (
            .O(N__33240),
            .I(N__33216));
    InMux I__6204 (
            .O(N__33239),
            .I(N__33213));
    InMux I__6203 (
            .O(N__33238),
            .I(N__33204));
    InMux I__6202 (
            .O(N__33237),
            .I(N__33204));
    InMux I__6201 (
            .O(N__33236),
            .I(N__33204));
    InMux I__6200 (
            .O(N__33235),
            .I(N__33204));
    InMux I__6199 (
            .O(N__33234),
            .I(N__33199));
    LocalMux I__6198 (
            .O(N__33231),
            .I(N__33196));
    InMux I__6197 (
            .O(N__33230),
            .I(N__33191));
    InMux I__6196 (
            .O(N__33229),
            .I(N__33191));
    InMux I__6195 (
            .O(N__33228),
            .I(N__33167));
    InMux I__6194 (
            .O(N__33227),
            .I(N__33167));
    InMux I__6193 (
            .O(N__33226),
            .I(N__33167));
    InMux I__6192 (
            .O(N__33225),
            .I(N__33167));
    InMux I__6191 (
            .O(N__33224),
            .I(N__33167));
    InMux I__6190 (
            .O(N__33223),
            .I(N__33167));
    LocalMux I__6189 (
            .O(N__33216),
            .I(N__33164));
    LocalMux I__6188 (
            .O(N__33213),
            .I(N__33159));
    LocalMux I__6187 (
            .O(N__33204),
            .I(N__33159));
    InMux I__6186 (
            .O(N__33203),
            .I(N__33154));
    InMux I__6185 (
            .O(N__33202),
            .I(N__33154));
    LocalMux I__6184 (
            .O(N__33199),
            .I(N__33151));
    Span4Mux_v I__6183 (
            .O(N__33196),
            .I(N__33146));
    LocalMux I__6182 (
            .O(N__33191),
            .I(N__33146));
    InMux I__6181 (
            .O(N__33190),
            .I(N__33135));
    InMux I__6180 (
            .O(N__33189),
            .I(N__33135));
    InMux I__6179 (
            .O(N__33188),
            .I(N__33135));
    InMux I__6178 (
            .O(N__33187),
            .I(N__33135));
    InMux I__6177 (
            .O(N__33186),
            .I(N__33135));
    InMux I__6176 (
            .O(N__33185),
            .I(N__33132));
    InMux I__6175 (
            .O(N__33184),
            .I(N__33127));
    InMux I__6174 (
            .O(N__33183),
            .I(N__33127));
    InMux I__6173 (
            .O(N__33182),
            .I(N__33122));
    InMux I__6172 (
            .O(N__33181),
            .I(N__33122));
    CascadeMux I__6171 (
            .O(N__33180),
            .I(N__33114));
    LocalMux I__6170 (
            .O(N__33167),
            .I(N__33107));
    Span4Mux_v I__6169 (
            .O(N__33164),
            .I(N__33107));
    Span4Mux_v I__6168 (
            .O(N__33159),
            .I(N__33107));
    LocalMux I__6167 (
            .O(N__33154),
            .I(N__33104));
    Span4Mux_v I__6166 (
            .O(N__33151),
            .I(N__33101));
    Span4Mux_h I__6165 (
            .O(N__33146),
            .I(N__33098));
    LocalMux I__6164 (
            .O(N__33135),
            .I(N__33095));
    LocalMux I__6163 (
            .O(N__33132),
            .I(N__33088));
    LocalMux I__6162 (
            .O(N__33127),
            .I(N__33088));
    LocalMux I__6161 (
            .O(N__33122),
            .I(N__33088));
    InMux I__6160 (
            .O(N__33121),
            .I(N__33085));
    InMux I__6159 (
            .O(N__33120),
            .I(N__33078));
    InMux I__6158 (
            .O(N__33119),
            .I(N__33078));
    InMux I__6157 (
            .O(N__33118),
            .I(N__33078));
    InMux I__6156 (
            .O(N__33117),
            .I(N__33073));
    InMux I__6155 (
            .O(N__33114),
            .I(N__33073));
    Sp12to4 I__6154 (
            .O(N__33107),
            .I(N__33070));
    Span4Mux_h I__6153 (
            .O(N__33104),
            .I(N__33067));
    Span4Mux_h I__6152 (
            .O(N__33101),
            .I(N__33062));
    Span4Mux_v I__6151 (
            .O(N__33098),
            .I(N__33062));
    Span4Mux_v I__6150 (
            .O(N__33095),
            .I(N__33057));
    Span4Mux_v I__6149 (
            .O(N__33088),
            .I(N__33057));
    LocalMux I__6148 (
            .O(N__33085),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    LocalMux I__6147 (
            .O(N__33078),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    LocalMux I__6146 (
            .O(N__33073),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    Odrv12 I__6145 (
            .O(N__33070),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    Odrv4 I__6144 (
            .O(N__33067),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    Odrv4 I__6143 (
            .O(N__33062),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    Odrv4 I__6142 (
            .O(N__33057),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    CascadeMux I__6141 (
            .O(N__33042),
            .I(N__33037));
    CascadeMux I__6140 (
            .O(N__33041),
            .I(N__33031));
    InMux I__6139 (
            .O(N__33040),
            .I(N__33026));
    InMux I__6138 (
            .O(N__33037),
            .I(N__33026));
    InMux I__6137 (
            .O(N__33036),
            .I(N__33023));
    InMux I__6136 (
            .O(N__33035),
            .I(N__33020));
    CascadeMux I__6135 (
            .O(N__33034),
            .I(N__33015));
    InMux I__6134 (
            .O(N__33031),
            .I(N__33012));
    LocalMux I__6133 (
            .O(N__33026),
            .I(N__33007));
    LocalMux I__6132 (
            .O(N__33023),
            .I(N__33007));
    LocalMux I__6131 (
            .O(N__33020),
            .I(N__33004));
    CascadeMux I__6130 (
            .O(N__33019),
            .I(N__33000));
    InMux I__6129 (
            .O(N__33018),
            .I(N__32992));
    InMux I__6128 (
            .O(N__33015),
            .I(N__32989));
    LocalMux I__6127 (
            .O(N__33012),
            .I(N__32986));
    Span4Mux_h I__6126 (
            .O(N__33007),
            .I(N__32983));
    Span4Mux_v I__6125 (
            .O(N__33004),
            .I(N__32980));
    InMux I__6124 (
            .O(N__33003),
            .I(N__32977));
    InMux I__6123 (
            .O(N__33000),
            .I(N__32974));
    InMux I__6122 (
            .O(N__32999),
            .I(N__32971));
    InMux I__6121 (
            .O(N__32998),
            .I(N__32968));
    InMux I__6120 (
            .O(N__32997),
            .I(N__32961));
    InMux I__6119 (
            .O(N__32996),
            .I(N__32961));
    InMux I__6118 (
            .O(N__32995),
            .I(N__32961));
    LocalMux I__6117 (
            .O(N__32992),
            .I(N__32958));
    LocalMux I__6116 (
            .O(N__32989),
            .I(N__32949));
    Span4Mux_v I__6115 (
            .O(N__32986),
            .I(N__32949));
    Span4Mux_v I__6114 (
            .O(N__32983),
            .I(N__32949));
    Span4Mux_h I__6113 (
            .O(N__32980),
            .I(N__32949));
    LocalMux I__6112 (
            .O(N__32977),
            .I(\phase_controller_inst1.stoper_hc.N_326 ));
    LocalMux I__6111 (
            .O(N__32974),
            .I(\phase_controller_inst1.stoper_hc.N_326 ));
    LocalMux I__6110 (
            .O(N__32971),
            .I(\phase_controller_inst1.stoper_hc.N_326 ));
    LocalMux I__6109 (
            .O(N__32968),
            .I(\phase_controller_inst1.stoper_hc.N_326 ));
    LocalMux I__6108 (
            .O(N__32961),
            .I(\phase_controller_inst1.stoper_hc.N_326 ));
    Odrv12 I__6107 (
            .O(N__32958),
            .I(\phase_controller_inst1.stoper_hc.N_326 ));
    Odrv4 I__6106 (
            .O(N__32949),
            .I(\phase_controller_inst1.stoper_hc.N_326 ));
    InMux I__6105 (
            .O(N__32934),
            .I(N__32931));
    LocalMux I__6104 (
            .O(N__32931),
            .I(N__32927));
    InMux I__6103 (
            .O(N__32930),
            .I(N__32924));
    Odrv4 I__6102 (
            .O(N__32927),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ));
    LocalMux I__6101 (
            .O(N__32924),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ));
    InMux I__6100 (
            .O(N__32919),
            .I(N__32916));
    LocalMux I__6099 (
            .O(N__32916),
            .I(N__32913));
    Span4Mux_v I__6098 (
            .O(N__32913),
            .I(N__32910));
    Span4Mux_h I__6097 (
            .O(N__32910),
            .I(N__32907));
    Span4Mux_v I__6096 (
            .O(N__32907),
            .I(N__32904));
    Odrv4 I__6095 (
            .O(N__32904),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CEMux I__6094 (
            .O(N__32901),
            .I(N__32893));
    CEMux I__6093 (
            .O(N__32900),
            .I(N__32890));
    CEMux I__6092 (
            .O(N__32899),
            .I(N__32886));
    CEMux I__6091 (
            .O(N__32898),
            .I(N__32883));
    CEMux I__6090 (
            .O(N__32897),
            .I(N__32880));
    CEMux I__6089 (
            .O(N__32896),
            .I(N__32876));
    LocalMux I__6088 (
            .O(N__32893),
            .I(N__32873));
    LocalMux I__6087 (
            .O(N__32890),
            .I(N__32870));
    CEMux I__6086 (
            .O(N__32889),
            .I(N__32867));
    LocalMux I__6085 (
            .O(N__32886),
            .I(N__32841));
    LocalMux I__6084 (
            .O(N__32883),
            .I(N__32838));
    LocalMux I__6083 (
            .O(N__32880),
            .I(N__32835));
    CEMux I__6082 (
            .O(N__32879),
            .I(N__32832));
    LocalMux I__6081 (
            .O(N__32876),
            .I(N__32827));
    Span4Mux_v I__6080 (
            .O(N__32873),
            .I(N__32827));
    Span4Mux_h I__6079 (
            .O(N__32870),
            .I(N__32824));
    LocalMux I__6078 (
            .O(N__32867),
            .I(N__32821));
    InMux I__6077 (
            .O(N__32866),
            .I(N__32812));
    InMux I__6076 (
            .O(N__32865),
            .I(N__32812));
    InMux I__6075 (
            .O(N__32864),
            .I(N__32812));
    InMux I__6074 (
            .O(N__32863),
            .I(N__32812));
    InMux I__6073 (
            .O(N__32862),
            .I(N__32803));
    InMux I__6072 (
            .O(N__32861),
            .I(N__32803));
    InMux I__6071 (
            .O(N__32860),
            .I(N__32803));
    InMux I__6070 (
            .O(N__32859),
            .I(N__32803));
    InMux I__6069 (
            .O(N__32858),
            .I(N__32794));
    InMux I__6068 (
            .O(N__32857),
            .I(N__32794));
    InMux I__6067 (
            .O(N__32856),
            .I(N__32794));
    InMux I__6066 (
            .O(N__32855),
            .I(N__32794));
    InMux I__6065 (
            .O(N__32854),
            .I(N__32785));
    InMux I__6064 (
            .O(N__32853),
            .I(N__32785));
    InMux I__6063 (
            .O(N__32852),
            .I(N__32785));
    InMux I__6062 (
            .O(N__32851),
            .I(N__32785));
    InMux I__6061 (
            .O(N__32850),
            .I(N__32778));
    InMux I__6060 (
            .O(N__32849),
            .I(N__32778));
    InMux I__6059 (
            .O(N__32848),
            .I(N__32778));
    InMux I__6058 (
            .O(N__32847),
            .I(N__32769));
    InMux I__6057 (
            .O(N__32846),
            .I(N__32769));
    InMux I__6056 (
            .O(N__32845),
            .I(N__32769));
    InMux I__6055 (
            .O(N__32844),
            .I(N__32769));
    Span4Mux_v I__6054 (
            .O(N__32841),
            .I(N__32766));
    Span4Mux_v I__6053 (
            .O(N__32838),
            .I(N__32751));
    Span4Mux_v I__6052 (
            .O(N__32835),
            .I(N__32751));
    LocalMux I__6051 (
            .O(N__32832),
            .I(N__32751));
    Span4Mux_h I__6050 (
            .O(N__32827),
            .I(N__32746));
    Span4Mux_v I__6049 (
            .O(N__32824),
            .I(N__32746));
    Span4Mux_v I__6048 (
            .O(N__32821),
            .I(N__32743));
    LocalMux I__6047 (
            .O(N__32812),
            .I(N__32730));
    LocalMux I__6046 (
            .O(N__32803),
            .I(N__32730));
    LocalMux I__6045 (
            .O(N__32794),
            .I(N__32730));
    LocalMux I__6044 (
            .O(N__32785),
            .I(N__32730));
    LocalMux I__6043 (
            .O(N__32778),
            .I(N__32730));
    LocalMux I__6042 (
            .O(N__32769),
            .I(N__32730));
    Span4Mux_v I__6041 (
            .O(N__32766),
            .I(N__32727));
    InMux I__6040 (
            .O(N__32765),
            .I(N__32724));
    InMux I__6039 (
            .O(N__32764),
            .I(N__32717));
    InMux I__6038 (
            .O(N__32763),
            .I(N__32717));
    InMux I__6037 (
            .O(N__32762),
            .I(N__32717));
    InMux I__6036 (
            .O(N__32761),
            .I(N__32708));
    InMux I__6035 (
            .O(N__32760),
            .I(N__32708));
    InMux I__6034 (
            .O(N__32759),
            .I(N__32708));
    InMux I__6033 (
            .O(N__32758),
            .I(N__32708));
    Span4Mux_v I__6032 (
            .O(N__32751),
            .I(N__32703));
    Span4Mux_v I__6031 (
            .O(N__32746),
            .I(N__32703));
    Span4Mux_h I__6030 (
            .O(N__32743),
            .I(N__32696));
    Span4Mux_v I__6029 (
            .O(N__32730),
            .I(N__32696));
    Span4Mux_h I__6028 (
            .O(N__32727),
            .I(N__32696));
    LocalMux I__6027 (
            .O(N__32724),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__6026 (
            .O(N__32717),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__6025 (
            .O(N__32708),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__6024 (
            .O(N__32703),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__6023 (
            .O(N__32696),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__6022 (
            .O(N__32685),
            .I(N__32682));
    LocalMux I__6021 (
            .O(N__32682),
            .I(N__32678));
    InMux I__6020 (
            .O(N__32681),
            .I(N__32675));
    Span4Mux_h I__6019 (
            .O(N__32678),
            .I(N__32670));
    LocalMux I__6018 (
            .O(N__32675),
            .I(N__32670));
    Span4Mux_h I__6017 (
            .O(N__32670),
            .I(N__32666));
    InMux I__6016 (
            .O(N__32669),
            .I(N__32663));
    Odrv4 I__6015 (
            .O(N__32666),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    LocalMux I__6014 (
            .O(N__32663),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__6013 (
            .O(N__32658),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__6012 (
            .O(N__32655),
            .I(N__32651));
    InMux I__6011 (
            .O(N__32654),
            .I(N__32647));
    LocalMux I__6010 (
            .O(N__32651),
            .I(N__32644));
    InMux I__6009 (
            .O(N__32650),
            .I(N__32641));
    LocalMux I__6008 (
            .O(N__32647),
            .I(N__32638));
    Span4Mux_h I__6007 (
            .O(N__32644),
            .I(N__32635));
    LocalMux I__6006 (
            .O(N__32641),
            .I(N__32632));
    Odrv12 I__6005 (
            .O(N__32638),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__6004 (
            .O(N__32635),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__6003 (
            .O(N__32632),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__6002 (
            .O(N__32625),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__6001 (
            .O(N__32622),
            .I(bfn_12_11_0_));
    InMux I__6000 (
            .O(N__32619),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__5999 (
            .O(N__32616),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    CascadeMux I__5998 (
            .O(N__32613),
            .I(N__32609));
    InMux I__5997 (
            .O(N__32612),
            .I(N__32606));
    InMux I__5996 (
            .O(N__32609),
            .I(N__32603));
    LocalMux I__5995 (
            .O(N__32606),
            .I(N__32600));
    LocalMux I__5994 (
            .O(N__32603),
            .I(N__32596));
    Span4Mux_v I__5993 (
            .O(N__32600),
            .I(N__32593));
    InMux I__5992 (
            .O(N__32599),
            .I(N__32590));
    Span4Mux_v I__5991 (
            .O(N__32596),
            .I(N__32587));
    Span4Mux_h I__5990 (
            .O(N__32593),
            .I(N__32582));
    LocalMux I__5989 (
            .O(N__32590),
            .I(N__32582));
    Odrv4 I__5988 (
            .O(N__32587),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__5987 (
            .O(N__32582),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__5986 (
            .O(N__32577),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__5985 (
            .O(N__32574),
            .I(N__32570));
    InMux I__5984 (
            .O(N__32573),
            .I(N__32567));
    LocalMux I__5983 (
            .O(N__32570),
            .I(N__32563));
    LocalMux I__5982 (
            .O(N__32567),
            .I(N__32560));
    InMux I__5981 (
            .O(N__32566),
            .I(N__32557));
    Span4Mux_h I__5980 (
            .O(N__32563),
            .I(N__32554));
    Span4Mux_h I__5979 (
            .O(N__32560),
            .I(N__32549));
    LocalMux I__5978 (
            .O(N__32557),
            .I(N__32549));
    Odrv4 I__5977 (
            .O(N__32554),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__5976 (
            .O(N__32549),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__5975 (
            .O(N__32544),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__5974 (
            .O(N__32541),
            .I(N__32536));
    InMux I__5973 (
            .O(N__32540),
            .I(N__32531));
    InMux I__5972 (
            .O(N__32539),
            .I(N__32531));
    LocalMux I__5971 (
            .O(N__32536),
            .I(N__32526));
    LocalMux I__5970 (
            .O(N__32531),
            .I(N__32526));
    Span4Mux_h I__5969 (
            .O(N__32526),
            .I(N__32523));
    Odrv4 I__5968 (
            .O(N__32523),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__5967 (
            .O(N__32520),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__5966 (
            .O(N__32517),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__5965 (
            .O(N__32514),
            .I(N__32511));
    LocalMux I__5964 (
            .O(N__32511),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ));
    InMux I__5963 (
            .O(N__32508),
            .I(N__32504));
    InMux I__5962 (
            .O(N__32507),
            .I(N__32500));
    LocalMux I__5961 (
            .O(N__32504),
            .I(N__32497));
    InMux I__5960 (
            .O(N__32503),
            .I(N__32494));
    LocalMux I__5959 (
            .O(N__32500),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    Odrv12 I__5958 (
            .O(N__32497),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    LocalMux I__5957 (
            .O(N__32494),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    InMux I__5956 (
            .O(N__32487),
            .I(N__32483));
    InMux I__5955 (
            .O(N__32486),
            .I(N__32480));
    LocalMux I__5954 (
            .O(N__32483),
            .I(N__32474));
    LocalMux I__5953 (
            .O(N__32480),
            .I(N__32474));
    InMux I__5952 (
            .O(N__32479),
            .I(N__32471));
    Odrv4 I__5951 (
            .O(N__32474),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    LocalMux I__5950 (
            .O(N__32471),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    InMux I__5949 (
            .O(N__32466),
            .I(N__32463));
    LocalMux I__5948 (
            .O(N__32463),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__5947 (
            .O(N__32460),
            .I(N__32457));
    LocalMux I__5946 (
            .O(N__32457),
            .I(N__32454));
    Span4Mux_h I__5945 (
            .O(N__32454),
            .I(N__32450));
    InMux I__5944 (
            .O(N__32453),
            .I(N__32447));
    Span4Mux_h I__5943 (
            .O(N__32450),
            .I(N__32442));
    LocalMux I__5942 (
            .O(N__32447),
            .I(N__32442));
    Odrv4 I__5941 (
            .O(N__32442),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__5940 (
            .O(N__32439),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__5939 (
            .O(N__32436),
            .I(N__32433));
    LocalMux I__5938 (
            .O(N__32433),
            .I(N__32430));
    Span4Mux_v I__5937 (
            .O(N__32430),
            .I(N__32426));
    InMux I__5936 (
            .O(N__32429),
            .I(N__32423));
    Span4Mux_h I__5935 (
            .O(N__32426),
            .I(N__32418));
    LocalMux I__5934 (
            .O(N__32423),
            .I(N__32418));
    Odrv4 I__5933 (
            .O(N__32418),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__5932 (
            .O(N__32415),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__5931 (
            .O(N__32412),
            .I(N__32409));
    LocalMux I__5930 (
            .O(N__32409),
            .I(N__32405));
    InMux I__5929 (
            .O(N__32408),
            .I(N__32402));
    Span12Mux_h I__5928 (
            .O(N__32405),
            .I(N__32399));
    LocalMux I__5927 (
            .O(N__32402),
            .I(N__32396));
    Odrv12 I__5926 (
            .O(N__32399),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv4 I__5925 (
            .O(N__32396),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__5924 (
            .O(N__32391),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__5923 (
            .O(N__32388),
            .I(N__32385));
    LocalMux I__5922 (
            .O(N__32385),
            .I(N__32380));
    InMux I__5921 (
            .O(N__32384),
            .I(N__32377));
    InMux I__5920 (
            .O(N__32383),
            .I(N__32374));
    Span4Mux_v I__5919 (
            .O(N__32380),
            .I(N__32367));
    LocalMux I__5918 (
            .O(N__32377),
            .I(N__32367));
    LocalMux I__5917 (
            .O(N__32374),
            .I(N__32367));
    Span4Mux_h I__5916 (
            .O(N__32367),
            .I(N__32364));
    Odrv4 I__5915 (
            .O(N__32364),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__5914 (
            .O(N__32361),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__5913 (
            .O(N__32358),
            .I(N__32355));
    LocalMux I__5912 (
            .O(N__32355),
            .I(N__32352));
    Span4Mux_h I__5911 (
            .O(N__32352),
            .I(N__32348));
    CascadeMux I__5910 (
            .O(N__32351),
            .I(N__32345));
    Span4Mux_h I__5909 (
            .O(N__32348),
            .I(N__32341));
    InMux I__5908 (
            .O(N__32345),
            .I(N__32336));
    InMux I__5907 (
            .O(N__32344),
            .I(N__32336));
    Odrv4 I__5906 (
            .O(N__32341),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    LocalMux I__5905 (
            .O(N__32336),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__5904 (
            .O(N__32331),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__5903 (
            .O(N__32328),
            .I(N__32323));
    InMux I__5902 (
            .O(N__32327),
            .I(N__32319));
    InMux I__5901 (
            .O(N__32326),
            .I(N__32316));
    LocalMux I__5900 (
            .O(N__32323),
            .I(N__32313));
    CascadeMux I__5899 (
            .O(N__32322),
            .I(N__32309));
    LocalMux I__5898 (
            .O(N__32319),
            .I(N__32306));
    LocalMux I__5897 (
            .O(N__32316),
            .I(N__32303));
    Span4Mux_v I__5896 (
            .O(N__32313),
            .I(N__32300));
    InMux I__5895 (
            .O(N__32312),
            .I(N__32295));
    InMux I__5894 (
            .O(N__32309),
            .I(N__32295));
    Span4Mux_v I__5893 (
            .O(N__32306),
            .I(N__32292));
    Odrv4 I__5892 (
            .O(N__32303),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__5891 (
            .O(N__32300),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__5890 (
            .O(N__32295),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__5889 (
            .O(N__32292),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__5888 (
            .O(N__32283),
            .I(N__32280));
    LocalMux I__5887 (
            .O(N__32280),
            .I(N__32277));
    Span4Mux_h I__5886 (
            .O(N__32277),
            .I(N__32274));
    Odrv4 I__5885 (
            .O(N__32274),
            .I(\current_shift_inst.PI_CTRL.integrator_i_17 ));
    CascadeMux I__5884 (
            .O(N__32271),
            .I(N__32267));
    InMux I__5883 (
            .O(N__32270),
            .I(N__32262));
    InMux I__5882 (
            .O(N__32267),
            .I(N__32259));
    CascadeMux I__5881 (
            .O(N__32266),
            .I(N__32255));
    InMux I__5880 (
            .O(N__32265),
            .I(N__32252));
    LocalMux I__5879 (
            .O(N__32262),
            .I(N__32249));
    LocalMux I__5878 (
            .O(N__32259),
            .I(N__32246));
    InMux I__5877 (
            .O(N__32258),
            .I(N__32241));
    InMux I__5876 (
            .O(N__32255),
            .I(N__32241));
    LocalMux I__5875 (
            .O(N__32252),
            .I(N__32238));
    Span4Mux_h I__5874 (
            .O(N__32249),
            .I(N__32233));
    Span4Mux_h I__5873 (
            .O(N__32246),
            .I(N__32233));
    LocalMux I__5872 (
            .O(N__32241),
            .I(N__32230));
    Span4Mux_h I__5871 (
            .O(N__32238),
            .I(N__32227));
    Odrv4 I__5870 (
            .O(N__32233),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv12 I__5869 (
            .O(N__32230),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__5868 (
            .O(N__32227),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__5867 (
            .O(N__32220),
            .I(N__32217));
    LocalMux I__5866 (
            .O(N__32217),
            .I(N__32214));
    Span4Mux_h I__5865 (
            .O(N__32214),
            .I(N__32211));
    Odrv4 I__5864 (
            .O(N__32211),
            .I(\current_shift_inst.PI_CTRL.integrator_i_18 ));
    CascadeMux I__5863 (
            .O(N__32208),
            .I(N__32205));
    InMux I__5862 (
            .O(N__32205),
            .I(N__32201));
    CascadeMux I__5861 (
            .O(N__32204),
            .I(N__32198));
    LocalMux I__5860 (
            .O(N__32201),
            .I(N__32194));
    InMux I__5859 (
            .O(N__32198),
            .I(N__32191));
    InMux I__5858 (
            .O(N__32197),
            .I(N__32188));
    Span4Mux_h I__5857 (
            .O(N__32194),
            .I(N__32185));
    LocalMux I__5856 (
            .O(N__32191),
            .I(N__32182));
    LocalMux I__5855 (
            .O(N__32188),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    Odrv4 I__5854 (
            .O(N__32185),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    Odrv4 I__5853 (
            .O(N__32182),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    CascadeMux I__5852 (
            .O(N__32175),
            .I(N__32172));
    InMux I__5851 (
            .O(N__32172),
            .I(N__32169));
    LocalMux I__5850 (
            .O(N__32169),
            .I(N__32164));
    InMux I__5849 (
            .O(N__32168),
            .I(N__32160));
    CascadeMux I__5848 (
            .O(N__32167),
            .I(N__32157));
    Span4Mux_h I__5847 (
            .O(N__32164),
            .I(N__32154));
    InMux I__5846 (
            .O(N__32163),
            .I(N__32150));
    LocalMux I__5845 (
            .O(N__32160),
            .I(N__32147));
    InMux I__5844 (
            .O(N__32157),
            .I(N__32144));
    Span4Mux_h I__5843 (
            .O(N__32154),
            .I(N__32141));
    InMux I__5842 (
            .O(N__32153),
            .I(N__32138));
    LocalMux I__5841 (
            .O(N__32150),
            .I(N__32135));
    Odrv4 I__5840 (
            .O(N__32147),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__5839 (
            .O(N__32144),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__5838 (
            .O(N__32141),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__5837 (
            .O(N__32138),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__5836 (
            .O(N__32135),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__5835 (
            .O(N__32124),
            .I(N__32121));
    LocalMux I__5834 (
            .O(N__32121),
            .I(N__32118));
    Span4Mux_v I__5833 (
            .O(N__32118),
            .I(N__32115));
    Odrv4 I__5832 (
            .O(N__32115),
            .I(\current_shift_inst.PI_CTRL.integrator_i_12 ));
    CascadeMux I__5831 (
            .O(N__32112),
            .I(N__32109));
    InMux I__5830 (
            .O(N__32109),
            .I(N__32105));
    InMux I__5829 (
            .O(N__32108),
            .I(N__32102));
    LocalMux I__5828 (
            .O(N__32105),
            .I(N__32099));
    LocalMux I__5827 (
            .O(N__32102),
            .I(N__32096));
    Span4Mux_v I__5826 (
            .O(N__32099),
            .I(N__32093));
    Span4Mux_v I__5825 (
            .O(N__32096),
            .I(N__32088));
    Span4Mux_h I__5824 (
            .O(N__32093),
            .I(N__32085));
    InMux I__5823 (
            .O(N__32092),
            .I(N__32080));
    InMux I__5822 (
            .O(N__32091),
            .I(N__32080));
    Odrv4 I__5821 (
            .O(N__32088),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__5820 (
            .O(N__32085),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__5819 (
            .O(N__32080),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__5818 (
            .O(N__32073),
            .I(N__32070));
    LocalMux I__5817 (
            .O(N__32070),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_5 ));
    CascadeMux I__5816 (
            .O(N__32067),
            .I(N__32064));
    InMux I__5815 (
            .O(N__32064),
            .I(N__32061));
    LocalMux I__5814 (
            .O(N__32061),
            .I(N__32058));
    Span4Mux_h I__5813 (
            .O(N__32058),
            .I(N__32055));
    Odrv4 I__5812 (
            .O(N__32055),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5 ));
    InMux I__5811 (
            .O(N__32052),
            .I(N__32049));
    LocalMux I__5810 (
            .O(N__32049),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    InMux I__5809 (
            .O(N__32046),
            .I(N__32043));
    LocalMux I__5808 (
            .O(N__32043),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ));
    InMux I__5807 (
            .O(N__32040),
            .I(N__32037));
    LocalMux I__5806 (
            .O(N__32037),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ));
    InMux I__5805 (
            .O(N__32034),
            .I(N__32031));
    LocalMux I__5804 (
            .O(N__32031),
            .I(N__32028));
    Glb2LocalMux I__5803 (
            .O(N__32028),
            .I(N__32025));
    GlobalMux I__5802 (
            .O(N__32025),
            .I(clk_12mhz));
    IoInMux I__5801 (
            .O(N__32022),
            .I(N__32019));
    LocalMux I__5800 (
            .O(N__32019),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    IoInMux I__5799 (
            .O(N__32016),
            .I(N__32013));
    LocalMux I__5798 (
            .O(N__32013),
            .I(N__32010));
    Span4Mux_s1_v I__5797 (
            .O(N__32010),
            .I(N__32007));
    Odrv4 I__5796 (
            .O(N__32007),
            .I(\delay_measurement_inst.delay_tr_timer.N_395_i ));
    ClkMux I__5795 (
            .O(N__32004),
            .I(N__32001));
    GlobalMux I__5794 (
            .O(N__32001),
            .I(N__31998));
    gio2CtrlBuf I__5793 (
            .O(N__31998),
            .I(delay_tr_input_c_g));
    InMux I__5792 (
            .O(N__31995),
            .I(N__31991));
    InMux I__5791 (
            .O(N__31994),
            .I(N__31988));
    LocalMux I__5790 (
            .O(N__31991),
            .I(N__31982));
    LocalMux I__5789 (
            .O(N__31988),
            .I(N__31982));
    InMux I__5788 (
            .O(N__31987),
            .I(N__31979));
    Span4Mux_v I__5787 (
            .O(N__31982),
            .I(N__31976));
    LocalMux I__5786 (
            .O(N__31979),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    Odrv4 I__5785 (
            .O(N__31976),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    InMux I__5784 (
            .O(N__31971),
            .I(N__31965));
    InMux I__5783 (
            .O(N__31970),
            .I(N__31962));
    InMux I__5782 (
            .O(N__31969),
            .I(N__31958));
    InMux I__5781 (
            .O(N__31968),
            .I(N__31955));
    LocalMux I__5780 (
            .O(N__31965),
            .I(N__31952));
    LocalMux I__5779 (
            .O(N__31962),
            .I(N__31949));
    InMux I__5778 (
            .O(N__31961),
            .I(N__31946));
    LocalMux I__5777 (
            .O(N__31958),
            .I(N__31941));
    LocalMux I__5776 (
            .O(N__31955),
            .I(N__31941));
    Span4Mux_h I__5775 (
            .O(N__31952),
            .I(N__31936));
    Span4Mux_v I__5774 (
            .O(N__31949),
            .I(N__31936));
    LocalMux I__5773 (
            .O(N__31946),
            .I(N__31933));
    Span4Mux_h I__5772 (
            .O(N__31941),
            .I(N__31930));
    Odrv4 I__5771 (
            .O(N__31936),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv12 I__5770 (
            .O(N__31933),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__5769 (
            .O(N__31930),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__5768 (
            .O(N__31923),
            .I(N__31920));
    LocalMux I__5767 (
            .O(N__31920),
            .I(N__31917));
    Span4Mux_v I__5766 (
            .O(N__31917),
            .I(N__31914));
    Span4Mux_h I__5765 (
            .O(N__31914),
            .I(N__31911));
    Odrv4 I__5764 (
            .O(N__31911),
            .I(\current_shift_inst.PI_CTRL.integrator_i_27 ));
    InMux I__5763 (
            .O(N__31908),
            .I(N__31904));
    CascadeMux I__5762 (
            .O(N__31907),
            .I(N__31901));
    LocalMux I__5761 (
            .O(N__31904),
            .I(N__31896));
    InMux I__5760 (
            .O(N__31901),
            .I(N__31893));
    InMux I__5759 (
            .O(N__31900),
            .I(N__31890));
    InMux I__5758 (
            .O(N__31899),
            .I(N__31887));
    Span4Mux_v I__5757 (
            .O(N__31896),
            .I(N__31881));
    LocalMux I__5756 (
            .O(N__31893),
            .I(N__31881));
    LocalMux I__5755 (
            .O(N__31890),
            .I(N__31878));
    LocalMux I__5754 (
            .O(N__31887),
            .I(N__31875));
    InMux I__5753 (
            .O(N__31886),
            .I(N__31872));
    Span4Mux_h I__5752 (
            .O(N__31881),
            .I(N__31867));
    Span4Mux_h I__5751 (
            .O(N__31878),
            .I(N__31867));
    Odrv4 I__5750 (
            .O(N__31875),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__5749 (
            .O(N__31872),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__5748 (
            .O(N__31867),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__5747 (
            .O(N__31860),
            .I(N__31857));
    LocalMux I__5746 (
            .O(N__31857),
            .I(N__31854));
    Span4Mux_h I__5745 (
            .O(N__31854),
            .I(N__31851));
    Odrv4 I__5744 (
            .O(N__31851),
            .I(\current_shift_inst.PI_CTRL.integrator_i_13 ));
    CascadeMux I__5743 (
            .O(N__31848),
            .I(N__31844));
    InMux I__5742 (
            .O(N__31847),
            .I(N__31840));
    InMux I__5741 (
            .O(N__31844),
            .I(N__31837));
    InMux I__5740 (
            .O(N__31843),
            .I(N__31832));
    LocalMux I__5739 (
            .O(N__31840),
            .I(N__31829));
    LocalMux I__5738 (
            .O(N__31837),
            .I(N__31826));
    InMux I__5737 (
            .O(N__31836),
            .I(N__31821));
    InMux I__5736 (
            .O(N__31835),
            .I(N__31821));
    LocalMux I__5735 (
            .O(N__31832),
            .I(N__31818));
    Span12Mux_h I__5734 (
            .O(N__31829),
            .I(N__31813));
    Span12Mux_s8_h I__5733 (
            .O(N__31826),
            .I(N__31813));
    LocalMux I__5732 (
            .O(N__31821),
            .I(N__31810));
    Span4Mux_h I__5731 (
            .O(N__31818),
            .I(N__31807));
    Odrv12 I__5730 (
            .O(N__31813),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv12 I__5729 (
            .O(N__31810),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__5728 (
            .O(N__31807),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__5727 (
            .O(N__31800),
            .I(N__31797));
    LocalMux I__5726 (
            .O(N__31797),
            .I(N__31794));
    Span4Mux_v I__5725 (
            .O(N__31794),
            .I(N__31791));
    Odrv4 I__5724 (
            .O(N__31791),
            .I(\current_shift_inst.PI_CTRL.integrator_i_22 ));
    InMux I__5723 (
            .O(N__31788),
            .I(N__31785));
    LocalMux I__5722 (
            .O(N__31785),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ));
    CascadeMux I__5721 (
            .O(N__31782),
            .I(N__31779));
    InMux I__5720 (
            .O(N__31779),
            .I(N__31776));
    LocalMux I__5719 (
            .O(N__31776),
            .I(N__31773));
    Span4Mux_h I__5718 (
            .O(N__31773),
            .I(N__31769));
    InMux I__5717 (
            .O(N__31772),
            .I(N__31766));
    Odrv4 I__5716 (
            .O(N__31769),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__5715 (
            .O(N__31766),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    CascadeMux I__5714 (
            .O(N__31761),
            .I(N__31757));
    InMux I__5713 (
            .O(N__31760),
            .I(N__31752));
    InMux I__5712 (
            .O(N__31757),
            .I(N__31752));
    LocalMux I__5711 (
            .O(N__31752),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    CascadeMux I__5710 (
            .O(N__31749),
            .I(N__31746));
    InMux I__5709 (
            .O(N__31746),
            .I(N__31743));
    LocalMux I__5708 (
            .O(N__31743),
            .I(N__31739));
    InMux I__5707 (
            .O(N__31742),
            .I(N__31736));
    Odrv12 I__5706 (
            .O(N__31739),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__5705 (
            .O(N__31736),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__5704 (
            .O(N__31731),
            .I(N__31728));
    LocalMux I__5703 (
            .O(N__31728),
            .I(N__31725));
    Odrv12 I__5702 (
            .O(N__31725),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19 ));
    CascadeMux I__5701 (
            .O(N__31722),
            .I(N__31719));
    InMux I__5700 (
            .O(N__31719),
            .I(N__31714));
    InMux I__5699 (
            .O(N__31718),
            .I(N__31711));
    InMux I__5698 (
            .O(N__31717),
            .I(N__31708));
    LocalMux I__5697 (
            .O(N__31714),
            .I(N__31701));
    LocalMux I__5696 (
            .O(N__31711),
            .I(N__31701));
    LocalMux I__5695 (
            .O(N__31708),
            .I(N__31698));
    InMux I__5694 (
            .O(N__31707),
            .I(N__31693));
    InMux I__5693 (
            .O(N__31706),
            .I(N__31693));
    Span4Mux_v I__5692 (
            .O(N__31701),
            .I(N__31686));
    Span4Mux_h I__5691 (
            .O(N__31698),
            .I(N__31686));
    LocalMux I__5690 (
            .O(N__31693),
            .I(N__31686));
    Odrv4 I__5689 (
            .O(N__31686),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__5688 (
            .O(N__31683),
            .I(N__31679));
    InMux I__5687 (
            .O(N__31682),
            .I(N__31676));
    LocalMux I__5686 (
            .O(N__31679),
            .I(N__31673));
    LocalMux I__5685 (
            .O(N__31676),
            .I(N__31670));
    Span12Mux_v I__5684 (
            .O(N__31673),
            .I(N__31667));
    Odrv12 I__5683 (
            .O(N__31670),
            .I(state_ns_i_a2_1));
    Odrv12 I__5682 (
            .O(N__31667),
            .I(state_ns_i_a2_1));
    InMux I__5681 (
            .O(N__31662),
            .I(N__31659));
    LocalMux I__5680 (
            .O(N__31659),
            .I(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ));
    InMux I__5679 (
            .O(N__31656),
            .I(N__31653));
    LocalMux I__5678 (
            .O(N__31653),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    CascadeMux I__5677 (
            .O(N__31650),
            .I(N__31645));
    InMux I__5676 (
            .O(N__31649),
            .I(N__31641));
    InMux I__5675 (
            .O(N__31648),
            .I(N__31638));
    InMux I__5674 (
            .O(N__31645),
            .I(N__31633));
    InMux I__5673 (
            .O(N__31644),
            .I(N__31633));
    LocalMux I__5672 (
            .O(N__31641),
            .I(N__31630));
    LocalMux I__5671 (
            .O(N__31638),
            .I(N__31627));
    LocalMux I__5670 (
            .O(N__31633),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__5669 (
            .O(N__31630),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__5668 (
            .O(N__31627),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    CascadeMux I__5667 (
            .O(N__31620),
            .I(N__31617));
    InMux I__5666 (
            .O(N__31617),
            .I(N__31614));
    LocalMux I__5665 (
            .O(N__31614),
            .I(N__31609));
    InMux I__5664 (
            .O(N__31613),
            .I(N__31606));
    InMux I__5663 (
            .O(N__31612),
            .I(N__31603));
    Span4Mux_v I__5662 (
            .O(N__31609),
            .I(N__31600));
    LocalMux I__5661 (
            .O(N__31606),
            .I(N__31597));
    LocalMux I__5660 (
            .O(N__31603),
            .I(N__31594));
    Span4Mux_h I__5659 (
            .O(N__31600),
            .I(N__31589));
    Span4Mux_h I__5658 (
            .O(N__31597),
            .I(N__31589));
    Span12Mux_h I__5657 (
            .O(N__31594),
            .I(N__31584));
    Sp12to4 I__5656 (
            .O(N__31589),
            .I(N__31584));
    Span12Mux_v I__5655 (
            .O(N__31584),
            .I(N__31581));
    Odrv12 I__5654 (
            .O(N__31581),
            .I(il_max_comp1_D2));
    CascadeMux I__5653 (
            .O(N__31578),
            .I(N__31574));
    InMux I__5652 (
            .O(N__31577),
            .I(N__31571));
    InMux I__5651 (
            .O(N__31574),
            .I(N__31568));
    LocalMux I__5650 (
            .O(N__31571),
            .I(N__31562));
    LocalMux I__5649 (
            .O(N__31568),
            .I(N__31562));
    InMux I__5648 (
            .O(N__31567),
            .I(N__31559));
    Span4Mux_v I__5647 (
            .O(N__31562),
            .I(N__31553));
    LocalMux I__5646 (
            .O(N__31559),
            .I(N__31553));
    InMux I__5645 (
            .O(N__31558),
            .I(N__31550));
    Span4Mux_h I__5644 (
            .O(N__31553),
            .I(N__31547));
    LocalMux I__5643 (
            .O(N__31550),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__5642 (
            .O(N__31547),
            .I(\phase_controller_inst1.hc_time_passed ));
    CascadeMux I__5641 (
            .O(N__31542),
            .I(N__31538));
    InMux I__5640 (
            .O(N__31541),
            .I(N__31534));
    InMux I__5639 (
            .O(N__31538),
            .I(N__31531));
    InMux I__5638 (
            .O(N__31537),
            .I(N__31528));
    LocalMux I__5637 (
            .O(N__31534),
            .I(N__31525));
    LocalMux I__5636 (
            .O(N__31531),
            .I(N__31521));
    LocalMux I__5635 (
            .O(N__31528),
            .I(N__31516));
    Span4Mux_v I__5634 (
            .O(N__31525),
            .I(N__31516));
    InMux I__5633 (
            .O(N__31524),
            .I(N__31513));
    Odrv4 I__5632 (
            .O(N__31521),
            .I(elapsed_time_ns_1_RNI5GT8E1_0_13));
    Odrv4 I__5631 (
            .O(N__31516),
            .I(elapsed_time_ns_1_RNI5GT8E1_0_13));
    LocalMux I__5630 (
            .O(N__31513),
            .I(elapsed_time_ns_1_RNI5GT8E1_0_13));
    CascadeMux I__5629 (
            .O(N__31506),
            .I(N__31499));
    CascadeMux I__5628 (
            .O(N__31505),
            .I(N__31496));
    CascadeMux I__5627 (
            .O(N__31504),
            .I(N__31490));
    InMux I__5626 (
            .O(N__31503),
            .I(N__31480));
    InMux I__5625 (
            .O(N__31502),
            .I(N__31480));
    InMux I__5624 (
            .O(N__31499),
            .I(N__31480));
    InMux I__5623 (
            .O(N__31496),
            .I(N__31480));
    InMux I__5622 (
            .O(N__31495),
            .I(N__31470));
    InMux I__5621 (
            .O(N__31494),
            .I(N__31470));
    InMux I__5620 (
            .O(N__31493),
            .I(N__31470));
    InMux I__5619 (
            .O(N__31490),
            .I(N__31470));
    InMux I__5618 (
            .O(N__31489),
            .I(N__31467));
    LocalMux I__5617 (
            .O(N__31480),
            .I(N__31464));
    InMux I__5616 (
            .O(N__31479),
            .I(N__31461));
    LocalMux I__5615 (
            .O(N__31470),
            .I(N__31456));
    LocalMux I__5614 (
            .O(N__31467),
            .I(N__31456));
    Span4Mux_v I__5613 (
            .O(N__31464),
            .I(N__31453));
    LocalMux I__5612 (
            .O(N__31461),
            .I(N__31448));
    Span4Mux_v I__5611 (
            .O(N__31456),
            .I(N__31448));
    Odrv4 I__5610 (
            .O(N__31453),
            .I(\phase_controller_inst1.stoper_hc.N_316 ));
    Odrv4 I__5609 (
            .O(N__31448),
            .I(\phase_controller_inst1.stoper_hc.N_316 ));
    CascadeMux I__5608 (
            .O(N__31443),
            .I(N__31434));
    CascadeMux I__5607 (
            .O(N__31442),
            .I(N__31426));
    CascadeMux I__5606 (
            .O(N__31441),
            .I(N__31422));
    CascadeMux I__5605 (
            .O(N__31440),
            .I(N__31419));
    InMux I__5604 (
            .O(N__31439),
            .I(N__31410));
    InMux I__5603 (
            .O(N__31438),
            .I(N__31410));
    InMux I__5602 (
            .O(N__31437),
            .I(N__31410));
    InMux I__5601 (
            .O(N__31434),
            .I(N__31410));
    InMux I__5600 (
            .O(N__31433),
            .I(N__31401));
    InMux I__5599 (
            .O(N__31432),
            .I(N__31401));
    InMux I__5598 (
            .O(N__31431),
            .I(N__31401));
    InMux I__5597 (
            .O(N__31430),
            .I(N__31401));
    InMux I__5596 (
            .O(N__31429),
            .I(N__31392));
    InMux I__5595 (
            .O(N__31426),
            .I(N__31389));
    InMux I__5594 (
            .O(N__31425),
            .I(N__31382));
    InMux I__5593 (
            .O(N__31422),
            .I(N__31382));
    InMux I__5592 (
            .O(N__31419),
            .I(N__31382));
    LocalMux I__5591 (
            .O(N__31410),
            .I(N__31377));
    LocalMux I__5590 (
            .O(N__31401),
            .I(N__31377));
    CascadeMux I__5589 (
            .O(N__31400),
            .I(N__31373));
    InMux I__5588 (
            .O(N__31399),
            .I(N__31359));
    InMux I__5587 (
            .O(N__31398),
            .I(N__31359));
    InMux I__5586 (
            .O(N__31397),
            .I(N__31359));
    InMux I__5585 (
            .O(N__31396),
            .I(N__31359));
    InMux I__5584 (
            .O(N__31395),
            .I(N__31359));
    LocalMux I__5583 (
            .O(N__31392),
            .I(N__31350));
    LocalMux I__5582 (
            .O(N__31389),
            .I(N__31350));
    LocalMux I__5581 (
            .O(N__31382),
            .I(N__31350));
    Span4Mux_v I__5580 (
            .O(N__31377),
            .I(N__31350));
    InMux I__5579 (
            .O(N__31376),
            .I(N__31347));
    InMux I__5578 (
            .O(N__31373),
            .I(N__31341));
    InMux I__5577 (
            .O(N__31372),
            .I(N__31334));
    InMux I__5576 (
            .O(N__31371),
            .I(N__31334));
    InMux I__5575 (
            .O(N__31370),
            .I(N__31334));
    LocalMux I__5574 (
            .O(N__31359),
            .I(N__31331));
    Span4Mux_v I__5573 (
            .O(N__31350),
            .I(N__31326));
    LocalMux I__5572 (
            .O(N__31347),
            .I(N__31326));
    InMux I__5571 (
            .O(N__31346),
            .I(N__31323));
    InMux I__5570 (
            .O(N__31345),
            .I(N__31318));
    InMux I__5569 (
            .O(N__31344),
            .I(N__31318));
    LocalMux I__5568 (
            .O(N__31341),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__5567 (
            .O(N__31334),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    Odrv4 I__5566 (
            .O(N__31331),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    Odrv4 I__5565 (
            .O(N__31326),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__5564 (
            .O(N__31323),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    LocalMux I__5563 (
            .O(N__31318),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    InMux I__5562 (
            .O(N__31305),
            .I(N__31301));
    InMux I__5561 (
            .O(N__31304),
            .I(N__31298));
    LocalMux I__5560 (
            .O(N__31301),
            .I(N__31295));
    LocalMux I__5559 (
            .O(N__31298),
            .I(N__31292));
    Span4Mux_v I__5558 (
            .O(N__31295),
            .I(N__31287));
    Span4Mux_h I__5557 (
            .O(N__31292),
            .I(N__31284));
    InMux I__5556 (
            .O(N__31291),
            .I(N__31279));
    InMux I__5555 (
            .O(N__31290),
            .I(N__31279));
    Odrv4 I__5554 (
            .O(N__31287),
            .I(elapsed_time_ns_1_RNIHHC6P1_0_18));
    Odrv4 I__5553 (
            .O(N__31284),
            .I(elapsed_time_ns_1_RNIHHC6P1_0_18));
    LocalMux I__5552 (
            .O(N__31279),
            .I(elapsed_time_ns_1_RNIHHC6P1_0_18));
    InMux I__5551 (
            .O(N__31272),
            .I(N__31269));
    LocalMux I__5550 (
            .O(N__31269),
            .I(N__31265));
    InMux I__5549 (
            .O(N__31268),
            .I(N__31262));
    Span4Mux_h I__5548 (
            .O(N__31265),
            .I(N__31259));
    LocalMux I__5547 (
            .O(N__31262),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    Odrv4 I__5546 (
            .O(N__31259),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__5545 (
            .O(N__31254),
            .I(N__31251));
    LocalMux I__5544 (
            .O(N__31251),
            .I(N__31248));
    Span4Mux_v I__5543 (
            .O(N__31248),
            .I(N__31244));
    InMux I__5542 (
            .O(N__31247),
            .I(N__31241));
    Odrv4 I__5541 (
            .O(N__31244),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    LocalMux I__5540 (
            .O(N__31241),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__5539 (
            .O(N__31236),
            .I(N__31232));
    InMux I__5538 (
            .O(N__31235),
            .I(N__31227));
    LocalMux I__5537 (
            .O(N__31232),
            .I(N__31224));
    InMux I__5536 (
            .O(N__31231),
            .I(N__31221));
    InMux I__5535 (
            .O(N__31230),
            .I(N__31218));
    LocalMux I__5534 (
            .O(N__31227),
            .I(N__31213));
    Span4Mux_v I__5533 (
            .O(N__31224),
            .I(N__31213));
    LocalMux I__5532 (
            .O(N__31221),
            .I(N__31210));
    LocalMux I__5531 (
            .O(N__31218),
            .I(elapsed_time_ns_1_RNIPKKEE1_0_8));
    Odrv4 I__5530 (
            .O(N__31213),
            .I(elapsed_time_ns_1_RNIPKKEE1_0_8));
    Odrv12 I__5529 (
            .O(N__31210),
            .I(elapsed_time_ns_1_RNIPKKEE1_0_8));
    InMux I__5528 (
            .O(N__31203),
            .I(N__31200));
    LocalMux I__5527 (
            .O(N__31200),
            .I(N__31196));
    InMux I__5526 (
            .O(N__31199),
            .I(N__31193));
    Odrv4 I__5525 (
            .O(N__31196),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__5524 (
            .O(N__31193),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__5523 (
            .O(N__31188),
            .I(N__31185));
    LocalMux I__5522 (
            .O(N__31185),
            .I(N__31181));
    InMux I__5521 (
            .O(N__31184),
            .I(N__31178));
    Odrv4 I__5520 (
            .O(N__31181),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    LocalMux I__5519 (
            .O(N__31178),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__5518 (
            .O(N__31173),
            .I(N__31169));
    CascadeMux I__5517 (
            .O(N__31172),
            .I(N__31166));
    LocalMux I__5516 (
            .O(N__31169),
            .I(N__31163));
    InMux I__5515 (
            .O(N__31166),
            .I(N__31160));
    Odrv4 I__5514 (
            .O(N__31163),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__5513 (
            .O(N__31160),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__5512 (
            .O(N__31155),
            .I(N__31152));
    LocalMux I__5511 (
            .O(N__31152),
            .I(N__31148));
    InMux I__5510 (
            .O(N__31151),
            .I(N__31145));
    Odrv4 I__5509 (
            .O(N__31148),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__5508 (
            .O(N__31145),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__5507 (
            .O(N__31140),
            .I(N__31137));
    LocalMux I__5506 (
            .O(N__31137),
            .I(N__31134));
    Sp12to4 I__5505 (
            .O(N__31134),
            .I(N__31131));
    Odrv12 I__5504 (
            .O(N__31131),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17 ));
    InMux I__5503 (
            .O(N__31128),
            .I(N__31125));
    LocalMux I__5502 (
            .O(N__31125),
            .I(N__31119));
    InMux I__5501 (
            .O(N__31124),
            .I(N__31116));
    InMux I__5500 (
            .O(N__31123),
            .I(N__31113));
    CascadeMux I__5499 (
            .O(N__31122),
            .I(N__31100));
    Span4Mux_v I__5498 (
            .O(N__31119),
            .I(N__31094));
    LocalMux I__5497 (
            .O(N__31116),
            .I(N__31094));
    LocalMux I__5496 (
            .O(N__31113),
            .I(N__31089));
    InMux I__5495 (
            .O(N__31112),
            .I(N__31086));
    CascadeMux I__5494 (
            .O(N__31111),
            .I(N__31082));
    CascadeMux I__5493 (
            .O(N__31110),
            .I(N__31077));
    CascadeMux I__5492 (
            .O(N__31109),
            .I(N__31074));
    CascadeMux I__5491 (
            .O(N__31108),
            .I(N__31069));
    CascadeMux I__5490 (
            .O(N__31107),
            .I(N__31063));
    InMux I__5489 (
            .O(N__31106),
            .I(N__31058));
    InMux I__5488 (
            .O(N__31105),
            .I(N__31058));
    CascadeMux I__5487 (
            .O(N__31104),
            .I(N__31052));
    InMux I__5486 (
            .O(N__31103),
            .I(N__31049));
    InMux I__5485 (
            .O(N__31100),
            .I(N__31044));
    InMux I__5484 (
            .O(N__31099),
            .I(N__31044));
    Span4Mux_v I__5483 (
            .O(N__31094),
            .I(N__31039));
    InMux I__5482 (
            .O(N__31093),
            .I(N__31036));
    InMux I__5481 (
            .O(N__31092),
            .I(N__31033));
    Span12Mux_h I__5480 (
            .O(N__31089),
            .I(N__31028));
    LocalMux I__5479 (
            .O(N__31086),
            .I(N__31028));
    InMux I__5478 (
            .O(N__31085),
            .I(N__31019));
    InMux I__5477 (
            .O(N__31082),
            .I(N__31019));
    InMux I__5476 (
            .O(N__31081),
            .I(N__31019));
    InMux I__5475 (
            .O(N__31080),
            .I(N__31019));
    InMux I__5474 (
            .O(N__31077),
            .I(N__31010));
    InMux I__5473 (
            .O(N__31074),
            .I(N__31010));
    InMux I__5472 (
            .O(N__31073),
            .I(N__31010));
    InMux I__5471 (
            .O(N__31072),
            .I(N__31010));
    InMux I__5470 (
            .O(N__31069),
            .I(N__30999));
    InMux I__5469 (
            .O(N__31068),
            .I(N__30999));
    InMux I__5468 (
            .O(N__31067),
            .I(N__30999));
    InMux I__5467 (
            .O(N__31066),
            .I(N__30999));
    InMux I__5466 (
            .O(N__31063),
            .I(N__30999));
    LocalMux I__5465 (
            .O(N__31058),
            .I(N__30996));
    InMux I__5464 (
            .O(N__31057),
            .I(N__30987));
    InMux I__5463 (
            .O(N__31056),
            .I(N__30987));
    InMux I__5462 (
            .O(N__31055),
            .I(N__30987));
    InMux I__5461 (
            .O(N__31052),
            .I(N__30987));
    LocalMux I__5460 (
            .O(N__31049),
            .I(N__30982));
    LocalMux I__5459 (
            .O(N__31044),
            .I(N__30982));
    InMux I__5458 (
            .O(N__31043),
            .I(N__30977));
    InMux I__5457 (
            .O(N__31042),
            .I(N__30977));
    Odrv4 I__5456 (
            .O(N__31039),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    LocalMux I__5455 (
            .O(N__31036),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    LocalMux I__5454 (
            .O(N__31033),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    Odrv12 I__5453 (
            .O(N__31028),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    LocalMux I__5452 (
            .O(N__31019),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    LocalMux I__5451 (
            .O(N__31010),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    LocalMux I__5450 (
            .O(N__30999),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    Odrv4 I__5449 (
            .O(N__30996),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    LocalMux I__5448 (
            .O(N__30987),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    Odrv4 I__5447 (
            .O(N__30982),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    LocalMux I__5446 (
            .O(N__30977),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk ));
    CascadeMux I__5445 (
            .O(N__30954),
            .I(N__30951));
    InMux I__5444 (
            .O(N__30951),
            .I(N__30946));
    InMux I__5443 (
            .O(N__30950),
            .I(N__30942));
    CascadeMux I__5442 (
            .O(N__30949),
            .I(N__30939));
    LocalMux I__5441 (
            .O(N__30946),
            .I(N__30935));
    InMux I__5440 (
            .O(N__30945),
            .I(N__30932));
    LocalMux I__5439 (
            .O(N__30942),
            .I(N__30929));
    InMux I__5438 (
            .O(N__30939),
            .I(N__30924));
    InMux I__5437 (
            .O(N__30938),
            .I(N__30924));
    Odrv4 I__5436 (
            .O(N__30935),
            .I(elapsed_time_ns_1_RNIIIC6P1_0_19));
    LocalMux I__5435 (
            .O(N__30932),
            .I(elapsed_time_ns_1_RNIIIC6P1_0_19));
    Odrv12 I__5434 (
            .O(N__30929),
            .I(elapsed_time_ns_1_RNIIIC6P1_0_19));
    LocalMux I__5433 (
            .O(N__30924),
            .I(elapsed_time_ns_1_RNIIIC6P1_0_19));
    InMux I__5432 (
            .O(N__30915),
            .I(N__30912));
    LocalMux I__5431 (
            .O(N__30912),
            .I(N__30909));
    Odrv4 I__5430 (
            .O(N__30909),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ));
    InMux I__5429 (
            .O(N__30906),
            .I(N__30903));
    LocalMux I__5428 (
            .O(N__30903),
            .I(N__30900));
    Span4Mux_v I__5427 (
            .O(N__30900),
            .I(N__30896));
    InMux I__5426 (
            .O(N__30899),
            .I(N__30893));
    Odrv4 I__5425 (
            .O(N__30896),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    LocalMux I__5424 (
            .O(N__30893),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    CascadeMux I__5423 (
            .O(N__30888),
            .I(N__30885));
    InMux I__5422 (
            .O(N__30885),
            .I(N__30882));
    LocalMux I__5421 (
            .O(N__30882),
            .I(N__30878));
    InMux I__5420 (
            .O(N__30881),
            .I(N__30875));
    Odrv12 I__5419 (
            .O(N__30878),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__5418 (
            .O(N__30875),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__5417 (
            .O(N__30870),
            .I(N__30866));
    CascadeMux I__5416 (
            .O(N__30869),
            .I(N__30863));
    LocalMux I__5415 (
            .O(N__30866),
            .I(N__30860));
    InMux I__5414 (
            .O(N__30863),
            .I(N__30857));
    Odrv12 I__5413 (
            .O(N__30860),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__5412 (
            .O(N__30857),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__5411 (
            .O(N__30852),
            .I(N__30849));
    LocalMux I__5410 (
            .O(N__30849),
            .I(N__30846));
    Span4Mux_v I__5409 (
            .O(N__30846),
            .I(N__30842));
    InMux I__5408 (
            .O(N__30845),
            .I(N__30839));
    Odrv4 I__5407 (
            .O(N__30842),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__5406 (
            .O(N__30839),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__5405 (
            .O(N__30834),
            .I(N__30831));
    LocalMux I__5404 (
            .O(N__30831),
            .I(N__30828));
    Odrv4 I__5403 (
            .O(N__30828),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18 ));
    InMux I__5402 (
            .O(N__30825),
            .I(N__30822));
    LocalMux I__5401 (
            .O(N__30822),
            .I(N__30818));
    InMux I__5400 (
            .O(N__30821),
            .I(N__30815));
    Odrv12 I__5399 (
            .O(N__30818),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    LocalMux I__5398 (
            .O(N__30815),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    CascadeMux I__5397 (
            .O(N__30810),
            .I(N__30807));
    InMux I__5396 (
            .O(N__30807),
            .I(N__30803));
    InMux I__5395 (
            .O(N__30806),
            .I(N__30800));
    LocalMux I__5394 (
            .O(N__30803),
            .I(N__30797));
    LocalMux I__5393 (
            .O(N__30800),
            .I(N__30794));
    Span4Mux_v I__5392 (
            .O(N__30797),
            .I(N__30791));
    Odrv4 I__5391 (
            .O(N__30794),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__5390 (
            .O(N__30791),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__5389 (
            .O(N__30786),
            .I(N__30782));
    InMux I__5388 (
            .O(N__30785),
            .I(N__30779));
    LocalMux I__5387 (
            .O(N__30782),
            .I(N__30776));
    LocalMux I__5386 (
            .O(N__30779),
            .I(N__30773));
    Span12Mux_v I__5385 (
            .O(N__30776),
            .I(N__30770));
    Span4Mux_h I__5384 (
            .O(N__30773),
            .I(N__30767));
    Odrv12 I__5383 (
            .O(N__30770),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__5382 (
            .O(N__30767),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__5381 (
            .O(N__30762),
            .I(N__30759));
    LocalMux I__5380 (
            .O(N__30759),
            .I(N__30755));
    InMux I__5379 (
            .O(N__30758),
            .I(N__30752));
    Span4Mux_h I__5378 (
            .O(N__30755),
            .I(N__30747));
    LocalMux I__5377 (
            .O(N__30752),
            .I(N__30747));
    Odrv4 I__5376 (
            .O(N__30747),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    CascadeMux I__5375 (
            .O(N__30744),
            .I(N__30740));
    InMux I__5374 (
            .O(N__30743),
            .I(N__30737));
    InMux I__5373 (
            .O(N__30740),
            .I(N__30734));
    LocalMux I__5372 (
            .O(N__30737),
            .I(N__30731));
    LocalMux I__5371 (
            .O(N__30734),
            .I(N__30728));
    Span4Mux_h I__5370 (
            .O(N__30731),
            .I(N__30723));
    Span4Mux_h I__5369 (
            .O(N__30728),
            .I(N__30723));
    Odrv4 I__5368 (
            .O(N__30723),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__5367 (
            .O(N__30720),
            .I(N__30717));
    LocalMux I__5366 (
            .O(N__30717),
            .I(N__30713));
    InMux I__5365 (
            .O(N__30716),
            .I(N__30710));
    Span4Mux_v I__5364 (
            .O(N__30713),
            .I(N__30707));
    LocalMux I__5363 (
            .O(N__30710),
            .I(N__30704));
    Odrv4 I__5362 (
            .O(N__30707),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__5361 (
            .O(N__30704),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    CascadeMux I__5360 (
            .O(N__30699),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16_cascade_ ));
    InMux I__5359 (
            .O(N__30696),
            .I(N__30693));
    LocalMux I__5358 (
            .O(N__30693),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25 ));
    CascadeMux I__5357 (
            .O(N__30690),
            .I(N__30687));
    InMux I__5356 (
            .O(N__30687),
            .I(N__30681));
    CascadeMux I__5355 (
            .O(N__30686),
            .I(N__30678));
    CascadeMux I__5354 (
            .O(N__30685),
            .I(N__30674));
    CascadeMux I__5353 (
            .O(N__30684),
            .I(N__30658));
    LocalMux I__5352 (
            .O(N__30681),
            .I(N__30652));
    InMux I__5351 (
            .O(N__30678),
            .I(N__30649));
    InMux I__5350 (
            .O(N__30677),
            .I(N__30644));
    InMux I__5349 (
            .O(N__30674),
            .I(N__30644));
    InMux I__5348 (
            .O(N__30673),
            .I(N__30641));
    InMux I__5347 (
            .O(N__30672),
            .I(N__30634));
    InMux I__5346 (
            .O(N__30671),
            .I(N__30634));
    InMux I__5345 (
            .O(N__30670),
            .I(N__30634));
    InMux I__5344 (
            .O(N__30669),
            .I(N__30627));
    InMux I__5343 (
            .O(N__30668),
            .I(N__30627));
    InMux I__5342 (
            .O(N__30667),
            .I(N__30627));
    InMux I__5341 (
            .O(N__30666),
            .I(N__30616));
    InMux I__5340 (
            .O(N__30665),
            .I(N__30616));
    InMux I__5339 (
            .O(N__30664),
            .I(N__30616));
    InMux I__5338 (
            .O(N__30663),
            .I(N__30616));
    InMux I__5337 (
            .O(N__30662),
            .I(N__30616));
    InMux I__5336 (
            .O(N__30661),
            .I(N__30607));
    InMux I__5335 (
            .O(N__30658),
            .I(N__30607));
    InMux I__5334 (
            .O(N__30657),
            .I(N__30607));
    InMux I__5333 (
            .O(N__30656),
            .I(N__30607));
    InMux I__5332 (
            .O(N__30655),
            .I(N__30604));
    Span4Mux_h I__5331 (
            .O(N__30652),
            .I(N__30597));
    LocalMux I__5330 (
            .O(N__30649),
            .I(N__30597));
    LocalMux I__5329 (
            .O(N__30644),
            .I(N__30597));
    LocalMux I__5328 (
            .O(N__30641),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    LocalMux I__5327 (
            .O(N__30634),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    LocalMux I__5326 (
            .O(N__30627),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    LocalMux I__5325 (
            .O(N__30616),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    LocalMux I__5324 (
            .O(N__30607),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    LocalMux I__5323 (
            .O(N__30604),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    Odrv4 I__5322 (
            .O(N__30597),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    InMux I__5321 (
            .O(N__30582),
            .I(N__30578));
    InMux I__5320 (
            .O(N__30581),
            .I(N__30575));
    LocalMux I__5319 (
            .O(N__30578),
            .I(elapsed_time_ns_1_RNI3FU8E1_0_20));
    LocalMux I__5318 (
            .O(N__30575),
            .I(elapsed_time_ns_1_RNI3FU8E1_0_20));
    CascadeMux I__5317 (
            .O(N__30570),
            .I(N__30567));
    InMux I__5316 (
            .O(N__30567),
            .I(N__30563));
    InMux I__5315 (
            .O(N__30566),
            .I(N__30559));
    LocalMux I__5314 (
            .O(N__30563),
            .I(N__30556));
    CascadeMux I__5313 (
            .O(N__30562),
            .I(N__30553));
    LocalMux I__5312 (
            .O(N__30559),
            .I(N__30548));
    Span4Mux_v I__5311 (
            .O(N__30556),
            .I(N__30548));
    InMux I__5310 (
            .O(N__30553),
            .I(N__30545));
    Odrv4 I__5309 (
            .O(N__30548),
            .I(elapsed_time_ns_1_RNI2DT8E1_0_10));
    LocalMux I__5308 (
            .O(N__30545),
            .I(elapsed_time_ns_1_RNI2DT8E1_0_10));
    CascadeMux I__5307 (
            .O(N__30540),
            .I(N__30535));
    InMux I__5306 (
            .O(N__30539),
            .I(N__30532));
    CascadeMux I__5305 (
            .O(N__30538),
            .I(N__30529));
    InMux I__5304 (
            .O(N__30535),
            .I(N__30526));
    LocalMux I__5303 (
            .O(N__30532),
            .I(N__30523));
    InMux I__5302 (
            .O(N__30529),
            .I(N__30519));
    LocalMux I__5301 (
            .O(N__30526),
            .I(N__30516));
    Span4Mux_v I__5300 (
            .O(N__30523),
            .I(N__30513));
    InMux I__5299 (
            .O(N__30522),
            .I(N__30510));
    LocalMux I__5298 (
            .O(N__30519),
            .I(elapsed_time_ns_1_RNI3ET8E1_0_11));
    Odrv12 I__5297 (
            .O(N__30516),
            .I(elapsed_time_ns_1_RNI3ET8E1_0_11));
    Odrv4 I__5296 (
            .O(N__30513),
            .I(elapsed_time_ns_1_RNI3ET8E1_0_11));
    LocalMux I__5295 (
            .O(N__30510),
            .I(elapsed_time_ns_1_RNI3ET8E1_0_11));
    CascadeMux I__5294 (
            .O(N__30501),
            .I(N__30498));
    InMux I__5293 (
            .O(N__30498),
            .I(N__30495));
    LocalMux I__5292 (
            .O(N__30495),
            .I(N__30490));
    InMux I__5291 (
            .O(N__30494),
            .I(N__30486));
    InMux I__5290 (
            .O(N__30493),
            .I(N__30483));
    Span4Mux_v I__5289 (
            .O(N__30490),
            .I(N__30480));
    InMux I__5288 (
            .O(N__30489),
            .I(N__30477));
    LocalMux I__5287 (
            .O(N__30486),
            .I(elapsed_time_ns_1_RNI4FT8E1_0_12));
    LocalMux I__5286 (
            .O(N__30483),
            .I(elapsed_time_ns_1_RNI4FT8E1_0_12));
    Odrv4 I__5285 (
            .O(N__30480),
            .I(elapsed_time_ns_1_RNI4FT8E1_0_12));
    LocalMux I__5284 (
            .O(N__30477),
            .I(elapsed_time_ns_1_RNI4FT8E1_0_12));
    InMux I__5283 (
            .O(N__30468),
            .I(N__30464));
    InMux I__5282 (
            .O(N__30467),
            .I(N__30461));
    LocalMux I__5281 (
            .O(N__30464),
            .I(elapsed_time_ns_1_RNI4GU8E1_0_21));
    LocalMux I__5280 (
            .O(N__30461),
            .I(elapsed_time_ns_1_RNI4GU8E1_0_21));
    CascadeMux I__5279 (
            .O(N__30456),
            .I(elapsed_time_ns_1_RNICOU8E1_0_29_cascade_));
    InMux I__5278 (
            .O(N__30453),
            .I(N__30450));
    LocalMux I__5277 (
            .O(N__30450),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15 ));
    CascadeMux I__5276 (
            .O(N__30447),
            .I(N__30444));
    InMux I__5275 (
            .O(N__30444),
            .I(N__30437));
    InMux I__5274 (
            .O(N__30443),
            .I(N__30437));
    InMux I__5273 (
            .O(N__30442),
            .I(N__30434));
    LocalMux I__5272 (
            .O(N__30437),
            .I(N__30429));
    LocalMux I__5271 (
            .O(N__30434),
            .I(N__30426));
    InMux I__5270 (
            .O(N__30433),
            .I(N__30423));
    InMux I__5269 (
            .O(N__30432),
            .I(N__30420));
    Span4Mux_v I__5268 (
            .O(N__30429),
            .I(N__30415));
    Span4Mux_h I__5267 (
            .O(N__30426),
            .I(N__30415));
    LocalMux I__5266 (
            .O(N__30423),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__5265 (
            .O(N__30420),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__5264 (
            .O(N__30415),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    InMux I__5263 (
            .O(N__30408),
            .I(N__30402));
    InMux I__5262 (
            .O(N__30407),
            .I(N__30402));
    LocalMux I__5261 (
            .O(N__30402),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__5260 (
            .O(N__30399),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__5259 (
            .O(N__30396),
            .I(N__30393));
    LocalMux I__5258 (
            .O(N__30393),
            .I(N__30386));
    InMux I__5257 (
            .O(N__30392),
            .I(N__30377));
    InMux I__5256 (
            .O(N__30391),
            .I(N__30377));
    InMux I__5255 (
            .O(N__30390),
            .I(N__30377));
    InMux I__5254 (
            .O(N__30389),
            .I(N__30377));
    Span4Mux_h I__5253 (
            .O(N__30386),
            .I(N__30374));
    LocalMux I__5252 (
            .O(N__30377),
            .I(N__30371));
    Odrv4 I__5251 (
            .O(N__30374),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv12 I__5250 (
            .O(N__30371),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    CascadeMux I__5249 (
            .O(N__30366),
            .I(N__30363));
    InMux I__5248 (
            .O(N__30363),
            .I(N__30359));
    InMux I__5247 (
            .O(N__30362),
            .I(N__30356));
    LocalMux I__5246 (
            .O(N__30359),
            .I(elapsed_time_ns_1_RNI8KU8E1_0_25));
    LocalMux I__5245 (
            .O(N__30356),
            .I(elapsed_time_ns_1_RNI8KU8E1_0_25));
    InMux I__5244 (
            .O(N__30351),
            .I(N__30347));
    InMux I__5243 (
            .O(N__30350),
            .I(N__30344));
    LocalMux I__5242 (
            .O(N__30347),
            .I(N__30339));
    LocalMux I__5241 (
            .O(N__30344),
            .I(N__30339));
    Span4Mux_v I__5240 (
            .O(N__30339),
            .I(N__30336));
    Odrv4 I__5239 (
            .O(N__30336),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    CascadeMux I__5238 (
            .O(N__30333),
            .I(elapsed_time_ns_1_RNI2DT8E1_0_10_cascade_));
    CascadeMux I__5237 (
            .O(N__30330),
            .I(N__30327));
    InMux I__5236 (
            .O(N__30327),
            .I(N__30324));
    LocalMux I__5235 (
            .O(N__30324),
            .I(N__30319));
    InMux I__5234 (
            .O(N__30323),
            .I(N__30316));
    InMux I__5233 (
            .O(N__30322),
            .I(N__30313));
    Span4Mux_h I__5232 (
            .O(N__30319),
            .I(N__30310));
    LocalMux I__5231 (
            .O(N__30316),
            .I(N__30305));
    LocalMux I__5230 (
            .O(N__30313),
            .I(N__30305));
    Odrv4 I__5229 (
            .O(N__30310),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ));
    Odrv4 I__5228 (
            .O(N__30305),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ));
    InMux I__5227 (
            .O(N__30300),
            .I(N__30297));
    LocalMux I__5226 (
            .O(N__30297),
            .I(N__30293));
    InMux I__5225 (
            .O(N__30296),
            .I(N__30290));
    Span4Mux_v I__5224 (
            .O(N__30293),
            .I(N__30287));
    LocalMux I__5223 (
            .O(N__30290),
            .I(N__30284));
    Odrv4 I__5222 (
            .O(N__30287),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv12 I__5221 (
            .O(N__30284),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__5220 (
            .O(N__30279),
            .I(N__30273));
    InMux I__5219 (
            .O(N__30278),
            .I(N__30273));
    LocalMux I__5218 (
            .O(N__30273),
            .I(elapsed_time_ns_1_RNI4HV8E1_0_30));
    InMux I__5217 (
            .O(N__30270),
            .I(N__30267));
    LocalMux I__5216 (
            .O(N__30267),
            .I(N__30264));
    Span4Mux_v I__5215 (
            .O(N__30264),
            .I(N__30261));
    Odrv4 I__5214 (
            .O(N__30261),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    CascadeMux I__5213 (
            .O(N__30258),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ));
    CascadeMux I__5212 (
            .O(N__30255),
            .I(N__30248));
    InMux I__5211 (
            .O(N__30254),
            .I(N__30245));
    InMux I__5210 (
            .O(N__30253),
            .I(N__30242));
    InMux I__5209 (
            .O(N__30252),
            .I(N__30239));
    InMux I__5208 (
            .O(N__30251),
            .I(N__30233));
    InMux I__5207 (
            .O(N__30248),
            .I(N__30233));
    LocalMux I__5206 (
            .O(N__30245),
            .I(N__30228));
    LocalMux I__5205 (
            .O(N__30242),
            .I(N__30225));
    LocalMux I__5204 (
            .O(N__30239),
            .I(N__30222));
    InMux I__5203 (
            .O(N__30238),
            .I(N__30219));
    LocalMux I__5202 (
            .O(N__30233),
            .I(N__30216));
    InMux I__5201 (
            .O(N__30232),
            .I(N__30213));
    InMux I__5200 (
            .O(N__30231),
            .I(N__30210));
    Odrv4 I__5199 (
            .O(N__30228),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    Odrv4 I__5198 (
            .O(N__30225),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    Odrv4 I__5197 (
            .O(N__30222),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    LocalMux I__5196 (
            .O(N__30219),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    Odrv4 I__5195 (
            .O(N__30216),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    LocalMux I__5194 (
            .O(N__30213),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    LocalMux I__5193 (
            .O(N__30210),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    InMux I__5192 (
            .O(N__30195),
            .I(N__30191));
    CascadeMux I__5191 (
            .O(N__30194),
            .I(N__30186));
    LocalMux I__5190 (
            .O(N__30191),
            .I(N__30183));
    InMux I__5189 (
            .O(N__30190),
            .I(N__30178));
    InMux I__5188 (
            .O(N__30189),
            .I(N__30178));
    InMux I__5187 (
            .O(N__30186),
            .I(N__30175));
    Span4Mux_h I__5186 (
            .O(N__30183),
            .I(N__30172));
    LocalMux I__5185 (
            .O(N__30178),
            .I(N__30169));
    LocalMux I__5184 (
            .O(N__30175),
            .I(elapsed_time_ns_1_RNIP93CP1_0_1));
    Odrv4 I__5183 (
            .O(N__30172),
            .I(elapsed_time_ns_1_RNIP93CP1_0_1));
    Odrv4 I__5182 (
            .O(N__30169),
            .I(elapsed_time_ns_1_RNIP93CP1_0_1));
    InMux I__5181 (
            .O(N__30162),
            .I(N__30159));
    LocalMux I__5180 (
            .O(N__30159),
            .I(N__30156));
    Span4Mux_v I__5179 (
            .O(N__30156),
            .I(N__30151));
    InMux I__5178 (
            .O(N__30155),
            .I(N__30144));
    InMux I__5177 (
            .O(N__30154),
            .I(N__30144));
    Span4Mux_h I__5176 (
            .O(N__30151),
            .I(N__30141));
    InMux I__5175 (
            .O(N__30150),
            .I(N__30136));
    InMux I__5174 (
            .O(N__30149),
            .I(N__30136));
    LocalMux I__5173 (
            .O(N__30144),
            .I(elapsed_time_ns_1_RNIRB3CP1_0_3));
    Odrv4 I__5172 (
            .O(N__30141),
            .I(elapsed_time_ns_1_RNIRB3CP1_0_3));
    LocalMux I__5171 (
            .O(N__30136),
            .I(elapsed_time_ns_1_RNIRB3CP1_0_3));
    CascadeMux I__5170 (
            .O(N__30129),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3_cascade_ ));
    InMux I__5169 (
            .O(N__30126),
            .I(N__30123));
    LocalMux I__5168 (
            .O(N__30123),
            .I(N__30119));
    InMux I__5167 (
            .O(N__30122),
            .I(N__30115));
    Span4Mux_v I__5166 (
            .O(N__30119),
            .I(N__30111));
    InMux I__5165 (
            .O(N__30118),
            .I(N__30108));
    LocalMux I__5164 (
            .O(N__30115),
            .I(N__30105));
    InMux I__5163 (
            .O(N__30114),
            .I(N__30102));
    Span4Mux_h I__5162 (
            .O(N__30111),
            .I(N__30099));
    LocalMux I__5161 (
            .O(N__30108),
            .I(N__30094));
    Span4Mux_h I__5160 (
            .O(N__30105),
            .I(N__30094));
    LocalMux I__5159 (
            .O(N__30102),
            .I(elapsed_time_ns_1_RNIOJKEE1_0_7));
    Odrv4 I__5158 (
            .O(N__30099),
            .I(elapsed_time_ns_1_RNIOJKEE1_0_7));
    Odrv4 I__5157 (
            .O(N__30094),
            .I(elapsed_time_ns_1_RNIOJKEE1_0_7));
    CascadeMux I__5156 (
            .O(N__30087),
            .I(N__30084));
    InMux I__5155 (
            .O(N__30084),
            .I(N__30079));
    InMux I__5154 (
            .O(N__30083),
            .I(N__30076));
    InMux I__5153 (
            .O(N__30082),
            .I(N__30073));
    LocalMux I__5152 (
            .O(N__30079),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ));
    LocalMux I__5151 (
            .O(N__30076),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ));
    LocalMux I__5150 (
            .O(N__30073),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ));
    CascadeMux I__5149 (
            .O(N__30066),
            .I(N__30059));
    InMux I__5148 (
            .O(N__30065),
            .I(N__30052));
    InMux I__5147 (
            .O(N__30064),
            .I(N__30052));
    InMux I__5146 (
            .O(N__30063),
            .I(N__30048));
    InMux I__5145 (
            .O(N__30062),
            .I(N__30045));
    InMux I__5144 (
            .O(N__30059),
            .I(N__30042));
    InMux I__5143 (
            .O(N__30058),
            .I(N__30039));
    InMux I__5142 (
            .O(N__30057),
            .I(N__30036));
    LocalMux I__5141 (
            .O(N__30052),
            .I(N__30033));
    InMux I__5140 (
            .O(N__30051),
            .I(N__30030));
    LocalMux I__5139 (
            .O(N__30048),
            .I(N__30027));
    LocalMux I__5138 (
            .O(N__30045),
            .I(N__30022));
    LocalMux I__5137 (
            .O(N__30042),
            .I(N__30022));
    LocalMux I__5136 (
            .O(N__30039),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15));
    LocalMux I__5135 (
            .O(N__30036),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15));
    Odrv4 I__5134 (
            .O(N__30033),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15));
    LocalMux I__5133 (
            .O(N__30030),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15));
    Odrv4 I__5132 (
            .O(N__30027),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15));
    Odrv4 I__5131 (
            .O(N__30022),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15));
    CascadeMux I__5130 (
            .O(N__30009),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ));
    CascadeMux I__5129 (
            .O(N__30006),
            .I(N__30002));
    InMux I__5128 (
            .O(N__30005),
            .I(N__29996));
    InMux I__5127 (
            .O(N__30002),
            .I(N__29996));
    InMux I__5126 (
            .O(N__30001),
            .I(N__29993));
    LocalMux I__5125 (
            .O(N__29996),
            .I(N__29990));
    LocalMux I__5124 (
            .O(N__29993),
            .I(elapsed_time_ns_1_RNIUE3CP1_0_6));
    Odrv4 I__5123 (
            .O(N__29990),
            .I(elapsed_time_ns_1_RNIUE3CP1_0_6));
    CascadeMux I__5122 (
            .O(N__29985),
            .I(\phase_controller_inst1.stoper_hc.N_328_cascade_ ));
    InMux I__5121 (
            .O(N__29982),
            .I(N__29978));
    CascadeMux I__5120 (
            .O(N__29981),
            .I(N__29975));
    LocalMux I__5119 (
            .O(N__29978),
            .I(N__29972));
    InMux I__5118 (
            .O(N__29975),
            .I(N__29969));
    Span4Mux_h I__5117 (
            .O(N__29972),
            .I(N__29966));
    LocalMux I__5116 (
            .O(N__29969),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    Odrv4 I__5115 (
            .O(N__29966),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    CascadeMux I__5114 (
            .O(N__29961),
            .I(N__29957));
    InMux I__5113 (
            .O(N__29960),
            .I(N__29952));
    InMux I__5112 (
            .O(N__29957),
            .I(N__29952));
    LocalMux I__5111 (
            .O(N__29952),
            .I(N__29947));
    InMux I__5110 (
            .O(N__29951),
            .I(N__29944));
    InMux I__5109 (
            .O(N__29950),
            .I(N__29941));
    Span4Mux_h I__5108 (
            .O(N__29947),
            .I(N__29938));
    LocalMux I__5107 (
            .O(N__29944),
            .I(N__29935));
    LocalMux I__5106 (
            .O(N__29941),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__5105 (
            .O(N__29938),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__5104 (
            .O(N__29935),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__5103 (
            .O(N__29928),
            .I(N__29925));
    LocalMux I__5102 (
            .O(N__29925),
            .I(N__29921));
    InMux I__5101 (
            .O(N__29924),
            .I(N__29918));
    Span4Mux_v I__5100 (
            .O(N__29921),
            .I(N__29915));
    LocalMux I__5099 (
            .O(N__29918),
            .I(N__29912));
    Odrv4 I__5098 (
            .O(N__29915),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    Odrv12 I__5097 (
            .O(N__29912),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__5096 (
            .O(N__29907),
            .I(N__29904));
    LocalMux I__5095 (
            .O(N__29904),
            .I(elapsed_time_ns_1_RNICOU8E1_0_29));
    InMux I__5094 (
            .O(N__29901),
            .I(N__29898));
    LocalMux I__5093 (
            .O(N__29898),
            .I(N__29895));
    Span4Mux_v I__5092 (
            .O(N__29895),
            .I(N__29892));
    Span4Mux_v I__5091 (
            .O(N__29892),
            .I(N__29889));
    Odrv4 I__5090 (
            .O(N__29889),
            .I(il_min_comp1_D1));
    InMux I__5089 (
            .O(N__29886),
            .I(N__29881));
    InMux I__5088 (
            .O(N__29885),
            .I(N__29876));
    InMux I__5087 (
            .O(N__29884),
            .I(N__29876));
    LocalMux I__5086 (
            .O(N__29881),
            .I(N__29871));
    LocalMux I__5085 (
            .O(N__29876),
            .I(N__29871));
    Odrv4 I__5084 (
            .O(N__29871),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ));
    InMux I__5083 (
            .O(N__29868),
            .I(N__29863));
    InMux I__5082 (
            .O(N__29867),
            .I(N__29860));
    InMux I__5081 (
            .O(N__29866),
            .I(N__29857));
    LocalMux I__5080 (
            .O(N__29863),
            .I(N__29854));
    LocalMux I__5079 (
            .O(N__29860),
            .I(N__29851));
    LocalMux I__5078 (
            .O(N__29857),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv4 I__5077 (
            .O(N__29854),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv4 I__5076 (
            .O(N__29851),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    InMux I__5075 (
            .O(N__29844),
            .I(N__29841));
    LocalMux I__5074 (
            .O(N__29841),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ));
    CascadeMux I__5073 (
            .O(N__29838),
            .I(N__29835));
    InMux I__5072 (
            .O(N__29835),
            .I(N__29832));
    LocalMux I__5071 (
            .O(N__29832),
            .I(N__29829));
    Odrv4 I__5070 (
            .O(N__29829),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0 ));
    InMux I__5069 (
            .O(N__29826),
            .I(N__29822));
    InMux I__5068 (
            .O(N__29825),
            .I(N__29819));
    LocalMux I__5067 (
            .O(N__29822),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    LocalMux I__5066 (
            .O(N__29819),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    InMux I__5065 (
            .O(N__29814),
            .I(N__29810));
    InMux I__5064 (
            .O(N__29813),
            .I(N__29807));
    LocalMux I__5063 (
            .O(N__29810),
            .I(N__29801));
    LocalMux I__5062 (
            .O(N__29807),
            .I(N__29798));
    InMux I__5061 (
            .O(N__29806),
            .I(N__29795));
    InMux I__5060 (
            .O(N__29805),
            .I(N__29792));
    InMux I__5059 (
            .O(N__29804),
            .I(N__29789));
    Span4Mux_v I__5058 (
            .O(N__29801),
            .I(N__29784));
    Span4Mux_v I__5057 (
            .O(N__29798),
            .I(N__29784));
    LocalMux I__5056 (
            .O(N__29795),
            .I(N__29779));
    LocalMux I__5055 (
            .O(N__29792),
            .I(N__29779));
    LocalMux I__5054 (
            .O(N__29789),
            .I(N__29776));
    Span4Mux_h I__5053 (
            .O(N__29784),
            .I(N__29773));
    Span4Mux_v I__5052 (
            .O(N__29779),
            .I(N__29770));
    Odrv12 I__5051 (
            .O(N__29776),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__5050 (
            .O(N__29773),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__5049 (
            .O(N__29770),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__5048 (
            .O(N__29763),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_ ));
    InMux I__5047 (
            .O(N__29760),
            .I(N__29757));
    LocalMux I__5046 (
            .O(N__29757),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ));
    CascadeMux I__5045 (
            .O(N__29754),
            .I(N__29751));
    InMux I__5044 (
            .O(N__29751),
            .I(N__29748));
    LocalMux I__5043 (
            .O(N__29748),
            .I(N__29745));
    Odrv12 I__5042 (
            .O(N__29745),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0 ));
    InMux I__5041 (
            .O(N__29742),
            .I(N__29738));
    CascadeMux I__5040 (
            .O(N__29741),
            .I(N__29735));
    LocalMux I__5039 (
            .O(N__29738),
            .I(N__29732));
    InMux I__5038 (
            .O(N__29735),
            .I(N__29729));
    Span4Mux_v I__5037 (
            .O(N__29732),
            .I(N__29726));
    LocalMux I__5036 (
            .O(N__29729),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__5035 (
            .O(N__29726),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__5034 (
            .O(N__29721),
            .I(N__29717));
    InMux I__5033 (
            .O(N__29720),
            .I(N__29714));
    LocalMux I__5032 (
            .O(N__29717),
            .I(N__29711));
    LocalMux I__5031 (
            .O(N__29714),
            .I(N__29708));
    Span4Mux_v I__5030 (
            .O(N__29711),
            .I(N__29703));
    Span4Mux_v I__5029 (
            .O(N__29708),
            .I(N__29703));
    Odrv4 I__5028 (
            .O(N__29703),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__5027 (
            .O(N__29700),
            .I(N__29697));
    LocalMux I__5026 (
            .O(N__29697),
            .I(N__29694));
    Span4Mux_h I__5025 (
            .O(N__29694),
            .I(N__29691));
    Odrv4 I__5024 (
            .O(N__29691),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15 ));
    InMux I__5023 (
            .O(N__29688),
            .I(N__29684));
    InMux I__5022 (
            .O(N__29687),
            .I(N__29681));
    LocalMux I__5021 (
            .O(N__29684),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2 ));
    LocalMux I__5020 (
            .O(N__29681),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2 ));
    CascadeMux I__5019 (
            .O(N__29676),
            .I(N__29673));
    InMux I__5018 (
            .O(N__29673),
            .I(N__29670));
    LocalMux I__5017 (
            .O(N__29670),
            .I(N__29667));
    Odrv4 I__5016 (
            .O(N__29667),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ));
    InMux I__5015 (
            .O(N__29664),
            .I(N__29660));
    InMux I__5014 (
            .O(N__29663),
            .I(N__29657));
    LocalMux I__5013 (
            .O(N__29660),
            .I(N__29652));
    LocalMux I__5012 (
            .O(N__29657),
            .I(N__29652));
    Span4Mux_h I__5011 (
            .O(N__29652),
            .I(N__29648));
    InMux I__5010 (
            .O(N__29651),
            .I(N__29645));
    Span4Mux_h I__5009 (
            .O(N__29648),
            .I(N__29642));
    LocalMux I__5008 (
            .O(N__29645),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    Odrv4 I__5007 (
            .O(N__29642),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    CascadeMux I__5006 (
            .O(N__29637),
            .I(N__29634));
    InMux I__5005 (
            .O(N__29634),
            .I(N__29631));
    LocalMux I__5004 (
            .O(N__29631),
            .I(N__29628));
    Sp12to4 I__5003 (
            .O(N__29628),
            .I(N__29625));
    Odrv12 I__5002 (
            .O(N__29625),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ));
    InMux I__5001 (
            .O(N__29622),
            .I(bfn_11_11_0_));
    InMux I__5000 (
            .O(N__29619),
            .I(N__29616));
    LocalMux I__4999 (
            .O(N__29616),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ));
    InMux I__4998 (
            .O(N__29613),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ));
    InMux I__4997 (
            .O(N__29610),
            .I(N__29606));
    InMux I__4996 (
            .O(N__29609),
            .I(N__29603));
    LocalMux I__4995 (
            .O(N__29606),
            .I(N__29598));
    LocalMux I__4994 (
            .O(N__29603),
            .I(N__29598));
    Span4Mux_h I__4993 (
            .O(N__29598),
            .I(N__29594));
    InMux I__4992 (
            .O(N__29597),
            .I(N__29591));
    Span4Mux_h I__4991 (
            .O(N__29594),
            .I(N__29588));
    LocalMux I__4990 (
            .O(N__29591),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv4 I__4989 (
            .O(N__29588),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    InMux I__4988 (
            .O(N__29583),
            .I(N__29580));
    LocalMux I__4987 (
            .O(N__29580),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ));
    InMux I__4986 (
            .O(N__29577),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ));
    InMux I__4985 (
            .O(N__29574),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ));
    InMux I__4984 (
            .O(N__29571),
            .I(N__29568));
    LocalMux I__4983 (
            .O(N__29568),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ));
    InMux I__4982 (
            .O(N__29565),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ));
    InMux I__4981 (
            .O(N__29562),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ));
    InMux I__4980 (
            .O(N__29559),
            .I(N__29556));
    LocalMux I__4979 (
            .O(N__29556),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ));
    InMux I__4978 (
            .O(N__29553),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ));
    InMux I__4977 (
            .O(N__29550),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_31 ));
    CascadeMux I__4976 (
            .O(N__29547),
            .I(N__29544));
    InMux I__4975 (
            .O(N__29544),
            .I(N__29541));
    LocalMux I__4974 (
            .O(N__29541),
            .I(N__29538));
    Span4Mux_h I__4973 (
            .O(N__29538),
            .I(N__29535));
    Odrv4 I__4972 (
            .O(N__29535),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0 ));
    CascadeMux I__4971 (
            .O(N__29532),
            .I(N__29529));
    InMux I__4970 (
            .O(N__29529),
            .I(N__29526));
    LocalMux I__4969 (
            .O(N__29526),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ));
    InMux I__4968 (
            .O(N__29523),
            .I(bfn_11_10_0_));
    InMux I__4967 (
            .O(N__29520),
            .I(N__29517));
    LocalMux I__4966 (
            .O(N__29517),
            .I(N__29512));
    InMux I__4965 (
            .O(N__29516),
            .I(N__29509));
    InMux I__4964 (
            .O(N__29515),
            .I(N__29506));
    Sp12to4 I__4963 (
            .O(N__29512),
            .I(N__29501));
    LocalMux I__4962 (
            .O(N__29509),
            .I(N__29501));
    LocalMux I__4961 (
            .O(N__29506),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    Odrv12 I__4960 (
            .O(N__29501),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    CascadeMux I__4959 (
            .O(N__29496),
            .I(N__29493));
    InMux I__4958 (
            .O(N__29493),
            .I(N__29490));
    LocalMux I__4957 (
            .O(N__29490),
            .I(N__29487));
    Odrv4 I__4956 (
            .O(N__29487),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ));
    InMux I__4955 (
            .O(N__29484),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ));
    CascadeMux I__4954 (
            .O(N__29481),
            .I(N__29478));
    InMux I__4953 (
            .O(N__29478),
            .I(N__29475));
    LocalMux I__4952 (
            .O(N__29475),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ));
    InMux I__4951 (
            .O(N__29472),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ));
    InMux I__4950 (
            .O(N__29469),
            .I(N__29466));
    LocalMux I__4949 (
            .O(N__29466),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ));
    InMux I__4948 (
            .O(N__29463),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ));
    InMux I__4947 (
            .O(N__29460),
            .I(N__29456));
    InMux I__4946 (
            .O(N__29459),
            .I(N__29453));
    LocalMux I__4945 (
            .O(N__29456),
            .I(N__29450));
    LocalMux I__4944 (
            .O(N__29453),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    Odrv4 I__4943 (
            .O(N__29450),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    InMux I__4942 (
            .O(N__29445),
            .I(N__29442));
    LocalMux I__4941 (
            .O(N__29442),
            .I(N__29439));
    Odrv4 I__4940 (
            .O(N__29439),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ));
    InMux I__4939 (
            .O(N__29436),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ));
    InMux I__4938 (
            .O(N__29433),
            .I(N__29430));
    LocalMux I__4937 (
            .O(N__29430),
            .I(N__29425));
    InMux I__4936 (
            .O(N__29429),
            .I(N__29422));
    InMux I__4935 (
            .O(N__29428),
            .I(N__29419));
    Span4Mux_v I__4934 (
            .O(N__29425),
            .I(N__29416));
    LocalMux I__4933 (
            .O(N__29422),
            .I(N__29413));
    LocalMux I__4932 (
            .O(N__29419),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv4 I__4931 (
            .O(N__29416),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv12 I__4930 (
            .O(N__29413),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    InMux I__4929 (
            .O(N__29406),
            .I(N__29403));
    LocalMux I__4928 (
            .O(N__29403),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ));
    InMux I__4927 (
            .O(N__29400),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ));
    InMux I__4926 (
            .O(N__29397),
            .I(N__29393));
    InMux I__4925 (
            .O(N__29396),
            .I(N__29390));
    LocalMux I__4924 (
            .O(N__29393),
            .I(N__29384));
    LocalMux I__4923 (
            .O(N__29390),
            .I(N__29384));
    InMux I__4922 (
            .O(N__29389),
            .I(N__29381));
    Span4Mux_v I__4921 (
            .O(N__29384),
            .I(N__29378));
    LocalMux I__4920 (
            .O(N__29381),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    Odrv4 I__4919 (
            .O(N__29378),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    InMux I__4918 (
            .O(N__29373),
            .I(N__29370));
    LocalMux I__4917 (
            .O(N__29370),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ));
    InMux I__4916 (
            .O(N__29367),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ));
    InMux I__4915 (
            .O(N__29364),
            .I(N__29359));
    InMux I__4914 (
            .O(N__29363),
            .I(N__29356));
    InMux I__4913 (
            .O(N__29362),
            .I(N__29353));
    LocalMux I__4912 (
            .O(N__29359),
            .I(N__29348));
    LocalMux I__4911 (
            .O(N__29356),
            .I(N__29348));
    LocalMux I__4910 (
            .O(N__29353),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    Odrv4 I__4909 (
            .O(N__29348),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    CascadeMux I__4908 (
            .O(N__29343),
            .I(N__29340));
    InMux I__4907 (
            .O(N__29340),
            .I(N__29337));
    LocalMux I__4906 (
            .O(N__29337),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ));
    InMux I__4905 (
            .O(N__29334),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ));
    InMux I__4904 (
            .O(N__29331),
            .I(N__29328));
    LocalMux I__4903 (
            .O(N__29328),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_8 ));
    InMux I__4902 (
            .O(N__29325),
            .I(bfn_11_9_0_));
    InMux I__4901 (
            .O(N__29322),
            .I(N__29319));
    LocalMux I__4900 (
            .O(N__29319),
            .I(N__29316));
    Span4Mux_h I__4899 (
            .O(N__29316),
            .I(N__29313));
    Odrv4 I__4898 (
            .O(N__29313),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_9 ));
    InMux I__4897 (
            .O(N__29310),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ));
    CascadeMux I__4896 (
            .O(N__29307),
            .I(N__29304));
    InMux I__4895 (
            .O(N__29304),
            .I(N__29301));
    LocalMux I__4894 (
            .O(N__29301),
            .I(N__29298));
    Odrv4 I__4893 (
            .O(N__29298),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_10 ));
    InMux I__4892 (
            .O(N__29295),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ));
    InMux I__4891 (
            .O(N__29292),
            .I(N__29289));
    LocalMux I__4890 (
            .O(N__29289),
            .I(N__29286));
    Odrv4 I__4889 (
            .O(N__29286),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_11 ));
    InMux I__4888 (
            .O(N__29283),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ));
    CascadeMux I__4887 (
            .O(N__29280),
            .I(N__29277));
    InMux I__4886 (
            .O(N__29277),
            .I(N__29274));
    LocalMux I__4885 (
            .O(N__29274),
            .I(N__29271));
    Odrv4 I__4884 (
            .O(N__29271),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_12 ));
    InMux I__4883 (
            .O(N__29268),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ));
    InMux I__4882 (
            .O(N__29265),
            .I(N__29262));
    LocalMux I__4881 (
            .O(N__29262),
            .I(N__29259));
    Span4Mux_h I__4880 (
            .O(N__29259),
            .I(N__29256));
    Odrv4 I__4879 (
            .O(N__29256),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    InMux I__4878 (
            .O(N__29253),
            .I(N__29250));
    LocalMux I__4877 (
            .O(N__29250),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_13 ));
    InMux I__4876 (
            .O(N__29247),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ));
    InMux I__4875 (
            .O(N__29244),
            .I(N__29241));
    LocalMux I__4874 (
            .O(N__29241),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ));
    InMux I__4873 (
            .O(N__29238),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ));
    CascadeMux I__4872 (
            .O(N__29235),
            .I(N__29232));
    InMux I__4871 (
            .O(N__29232),
            .I(N__29229));
    LocalMux I__4870 (
            .O(N__29229),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ));
    InMux I__4869 (
            .O(N__29226),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ));
    CascadeMux I__4868 (
            .O(N__29223),
            .I(N__29218));
    InMux I__4867 (
            .O(N__29222),
            .I(N__29215));
    CascadeMux I__4866 (
            .O(N__29221),
            .I(N__29211));
    InMux I__4865 (
            .O(N__29218),
            .I(N__29208));
    LocalMux I__4864 (
            .O(N__29215),
            .I(N__29205));
    InMux I__4863 (
            .O(N__29214),
            .I(N__29202));
    InMux I__4862 (
            .O(N__29211),
            .I(N__29199));
    LocalMux I__4861 (
            .O(N__29208),
            .I(N__29196));
    Span4Mux_h I__4860 (
            .O(N__29205),
            .I(N__29193));
    LocalMux I__4859 (
            .O(N__29202),
            .I(N__29190));
    LocalMux I__4858 (
            .O(N__29199),
            .I(N__29187));
    Span4Mux_h I__4857 (
            .O(N__29196),
            .I(N__29184));
    Span4Mux_v I__4856 (
            .O(N__29193),
            .I(N__29181));
    Span4Mux_v I__4855 (
            .O(N__29190),
            .I(N__29176));
    Span4Mux_h I__4854 (
            .O(N__29187),
            .I(N__29176));
    Odrv4 I__4853 (
            .O(N__29184),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__4852 (
            .O(N__29181),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__4851 (
            .O(N__29176),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    CascadeMux I__4850 (
            .O(N__29169),
            .I(N__29166));
    InMux I__4849 (
            .O(N__29166),
            .I(N__29163));
    LocalMux I__4848 (
            .O(N__29163),
            .I(N__29160));
    Span12Mux_v I__4847 (
            .O(N__29160),
            .I(N__29157));
    Odrv12 I__4846 (
            .O(N__29157),
            .I(\current_shift_inst.PI_CTRL.integrator_i_28 ));
    InMux I__4845 (
            .O(N__29154),
            .I(N__29151));
    LocalMux I__4844 (
            .O(N__29151),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ));
    InMux I__4843 (
            .O(N__29148),
            .I(N__29145));
    LocalMux I__4842 (
            .O(N__29145),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ));
    InMux I__4841 (
            .O(N__29142),
            .I(N__29139));
    LocalMux I__4840 (
            .O(N__29139),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ));
    InMux I__4839 (
            .O(N__29136),
            .I(N__29133));
    LocalMux I__4838 (
            .O(N__29133),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ));
    InMux I__4837 (
            .O(N__29130),
            .I(N__29127));
    LocalMux I__4836 (
            .O(N__29127),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ));
    InMux I__4835 (
            .O(N__29124),
            .I(N__29121));
    LocalMux I__4834 (
            .O(N__29121),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_4 ));
    InMux I__4833 (
            .O(N__29118),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ));
    InMux I__4832 (
            .O(N__29115),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ));
    InMux I__4831 (
            .O(N__29112),
            .I(N__29109));
    LocalMux I__4830 (
            .O(N__29109),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_6 ));
    InMux I__4829 (
            .O(N__29106),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ));
    InMux I__4828 (
            .O(N__29103),
            .I(N__29100));
    LocalMux I__4827 (
            .O(N__29100),
            .I(N__29097));
    Odrv4 I__4826 (
            .O(N__29097),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_7 ));
    InMux I__4825 (
            .O(N__29094),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ));
    CascadeMux I__4824 (
            .O(N__29091),
            .I(N__29087));
    InMux I__4823 (
            .O(N__29090),
            .I(N__29084));
    InMux I__4822 (
            .O(N__29087),
            .I(N__29080));
    LocalMux I__4821 (
            .O(N__29084),
            .I(N__29077));
    InMux I__4820 (
            .O(N__29083),
            .I(N__29074));
    LocalMux I__4819 (
            .O(N__29080),
            .I(N__29071));
    Span4Mux_v I__4818 (
            .O(N__29077),
            .I(N__29066));
    LocalMux I__4817 (
            .O(N__29074),
            .I(N__29066));
    Span4Mux_v I__4816 (
            .O(N__29071),
            .I(N__29061));
    Span4Mux_v I__4815 (
            .O(N__29066),
            .I(N__29058));
    InMux I__4814 (
            .O(N__29065),
            .I(N__29053));
    InMux I__4813 (
            .O(N__29064),
            .I(N__29053));
    Odrv4 I__4812 (
            .O(N__29061),
            .I(elapsed_time_ns_1_RNIGGC6P1_0_17));
    Odrv4 I__4811 (
            .O(N__29058),
            .I(elapsed_time_ns_1_RNIGGC6P1_0_17));
    LocalMux I__4810 (
            .O(N__29053),
            .I(elapsed_time_ns_1_RNIGGC6P1_0_17));
    CascadeMux I__4809 (
            .O(N__29046),
            .I(N__29042));
    InMux I__4808 (
            .O(N__29045),
            .I(N__29037));
    InMux I__4807 (
            .O(N__29042),
            .I(N__29037));
    LocalMux I__4806 (
            .O(N__29037),
            .I(N__29034));
    Odrv4 I__4805 (
            .O(N__29034),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__4804 (
            .O(N__29031),
            .I(N__29028));
    LocalMux I__4803 (
            .O(N__29028),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__4802 (
            .O(N__29025),
            .I(N__29021));
    InMux I__4801 (
            .O(N__29024),
            .I(N__29016));
    InMux I__4800 (
            .O(N__29021),
            .I(N__29016));
    LocalMux I__4799 (
            .O(N__29016),
            .I(N__29013));
    Odrv4 I__4798 (
            .O(N__29013),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__4797 (
            .O(N__29010),
            .I(N__29007));
    LocalMux I__4796 (
            .O(N__29007),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__4795 (
            .O(N__29004),
            .I(N__29000));
    CascadeMux I__4794 (
            .O(N__29003),
            .I(N__28994));
    InMux I__4793 (
            .O(N__29000),
            .I(N__28991));
    InMux I__4792 (
            .O(N__28999),
            .I(N__28988));
    InMux I__4791 (
            .O(N__28998),
            .I(N__28985));
    InMux I__4790 (
            .O(N__28997),
            .I(N__28982));
    InMux I__4789 (
            .O(N__28994),
            .I(N__28979));
    LocalMux I__4788 (
            .O(N__28991),
            .I(N__28976));
    LocalMux I__4787 (
            .O(N__28988),
            .I(N__28973));
    LocalMux I__4786 (
            .O(N__28985),
            .I(N__28970));
    LocalMux I__4785 (
            .O(N__28982),
            .I(N__28967));
    LocalMux I__4784 (
            .O(N__28979),
            .I(N__28962));
    Span4Mux_h I__4783 (
            .O(N__28976),
            .I(N__28962));
    Span4Mux_h I__4782 (
            .O(N__28973),
            .I(N__28957));
    Span4Mux_h I__4781 (
            .O(N__28970),
            .I(N__28957));
    Odrv4 I__4780 (
            .O(N__28967),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__4779 (
            .O(N__28962),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__4778 (
            .O(N__28957),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__4777 (
            .O(N__28950),
            .I(N__28947));
    LocalMux I__4776 (
            .O(N__28947),
            .I(N__28944));
    Span4Mux_h I__4775 (
            .O(N__28944),
            .I(N__28941));
    Odrv4 I__4774 (
            .O(N__28941),
            .I(\current_shift_inst.PI_CTRL.integrator_i_14 ));
    InMux I__4773 (
            .O(N__28938),
            .I(N__28934));
    InMux I__4772 (
            .O(N__28937),
            .I(N__28930));
    LocalMux I__4771 (
            .O(N__28934),
            .I(N__28926));
    InMux I__4770 (
            .O(N__28933),
            .I(N__28923));
    LocalMux I__4769 (
            .O(N__28930),
            .I(N__28920));
    InMux I__4768 (
            .O(N__28929),
            .I(N__28917));
    Span4Mux_h I__4767 (
            .O(N__28926),
            .I(N__28914));
    LocalMux I__4766 (
            .O(N__28923),
            .I(N__28911));
    Odrv4 I__4765 (
            .O(N__28920),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__4764 (
            .O(N__28917),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__4763 (
            .O(N__28914),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv12 I__4762 (
            .O(N__28911),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__4761 (
            .O(N__28902),
            .I(N__28899));
    LocalMux I__4760 (
            .O(N__28899),
            .I(N__28896));
    Span4Mux_h I__4759 (
            .O(N__28896),
            .I(N__28893));
    Odrv4 I__4758 (
            .O(N__28893),
            .I(\current_shift_inst.PI_CTRL.integrator_i_2 ));
    InMux I__4757 (
            .O(N__28890),
            .I(N__28884));
    InMux I__4756 (
            .O(N__28889),
            .I(N__28884));
    LocalMux I__4755 (
            .O(N__28884),
            .I(N__28880));
    InMux I__4754 (
            .O(N__28883),
            .I(N__28877));
    Span4Mux_v I__4753 (
            .O(N__28880),
            .I(N__28874));
    LocalMux I__4752 (
            .O(N__28877),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__4751 (
            .O(N__28874),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__4750 (
            .O(N__28869),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__4749 (
            .O(N__28866),
            .I(N__28860));
    InMux I__4748 (
            .O(N__28865),
            .I(N__28860));
    LocalMux I__4747 (
            .O(N__28860),
            .I(N__28856));
    InMux I__4746 (
            .O(N__28859),
            .I(N__28853));
    Span4Mux_v I__4745 (
            .O(N__28856),
            .I(N__28850));
    LocalMux I__4744 (
            .O(N__28853),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__4743 (
            .O(N__28850),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__4742 (
            .O(N__28845),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__4741 (
            .O(N__28842),
            .I(N__28838));
    CascadeMux I__4740 (
            .O(N__28841),
            .I(N__28835));
    InMux I__4739 (
            .O(N__28838),
            .I(N__28832));
    InMux I__4738 (
            .O(N__28835),
            .I(N__28829));
    LocalMux I__4737 (
            .O(N__28832),
            .I(N__28823));
    LocalMux I__4736 (
            .O(N__28829),
            .I(N__28823));
    InMux I__4735 (
            .O(N__28828),
            .I(N__28820));
    Span4Mux_v I__4734 (
            .O(N__28823),
            .I(N__28817));
    LocalMux I__4733 (
            .O(N__28820),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__4732 (
            .O(N__28817),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    CascadeMux I__4731 (
            .O(N__28812),
            .I(N__28808));
    InMux I__4730 (
            .O(N__28811),
            .I(N__28803));
    InMux I__4729 (
            .O(N__28808),
            .I(N__28803));
    LocalMux I__4728 (
            .O(N__28803),
            .I(N__28800));
    Odrv12 I__4727 (
            .O(N__28800),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__4726 (
            .O(N__28797),
            .I(bfn_10_22_0_));
    CascadeMux I__4725 (
            .O(N__28794),
            .I(N__28790));
    CascadeMux I__4724 (
            .O(N__28793),
            .I(N__28787));
    InMux I__4723 (
            .O(N__28790),
            .I(N__28784));
    InMux I__4722 (
            .O(N__28787),
            .I(N__28781));
    LocalMux I__4721 (
            .O(N__28784),
            .I(N__28776));
    LocalMux I__4720 (
            .O(N__28781),
            .I(N__28776));
    Span4Mux_v I__4719 (
            .O(N__28776),
            .I(N__28772));
    InMux I__4718 (
            .O(N__28775),
            .I(N__28769));
    Span4Mux_h I__4717 (
            .O(N__28772),
            .I(N__28766));
    LocalMux I__4716 (
            .O(N__28769),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__4715 (
            .O(N__28766),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__4714 (
            .O(N__28761),
            .I(N__28757));
    InMux I__4713 (
            .O(N__28760),
            .I(N__28754));
    LocalMux I__4712 (
            .O(N__28757),
            .I(N__28751));
    LocalMux I__4711 (
            .O(N__28754),
            .I(N__28748));
    Span4Mux_v I__4710 (
            .O(N__28751),
            .I(N__28743));
    Span4Mux_v I__4709 (
            .O(N__28748),
            .I(N__28743));
    Odrv4 I__4708 (
            .O(N__28743),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__4707 (
            .O(N__28740),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__4706 (
            .O(N__28737),
            .I(N__28730));
    InMux I__4705 (
            .O(N__28736),
            .I(N__28730));
    InMux I__4704 (
            .O(N__28735),
            .I(N__28727));
    LocalMux I__4703 (
            .O(N__28730),
            .I(N__28724));
    LocalMux I__4702 (
            .O(N__28727),
            .I(N__28719));
    Span4Mux_v I__4701 (
            .O(N__28724),
            .I(N__28719));
    Odrv4 I__4700 (
            .O(N__28719),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    CascadeMux I__4699 (
            .O(N__28716),
            .I(N__28713));
    InMux I__4698 (
            .O(N__28713),
            .I(N__28710));
    LocalMux I__4697 (
            .O(N__28710),
            .I(N__28706));
    InMux I__4696 (
            .O(N__28709),
            .I(N__28703));
    Span4Mux_v I__4695 (
            .O(N__28706),
            .I(N__28700));
    LocalMux I__4694 (
            .O(N__28703),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv4 I__4693 (
            .O(N__28700),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__4692 (
            .O(N__28695),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__4691 (
            .O(N__28692),
            .I(N__28689));
    LocalMux I__4690 (
            .O(N__28689),
            .I(N__28685));
    InMux I__4689 (
            .O(N__28688),
            .I(N__28682));
    Span4Mux_v I__4688 (
            .O(N__28685),
            .I(N__28679));
    LocalMux I__4687 (
            .O(N__28682),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv4 I__4686 (
            .O(N__28679),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__4685 (
            .O(N__28674),
            .I(N__28671));
    InMux I__4684 (
            .O(N__28671),
            .I(N__28667));
    InMux I__4683 (
            .O(N__28670),
            .I(N__28664));
    LocalMux I__4682 (
            .O(N__28667),
            .I(N__28659));
    LocalMux I__4681 (
            .O(N__28664),
            .I(N__28659));
    Span4Mux_h I__4680 (
            .O(N__28659),
            .I(N__28655));
    InMux I__4679 (
            .O(N__28658),
            .I(N__28652));
    Span4Mux_v I__4678 (
            .O(N__28655),
            .I(N__28649));
    LocalMux I__4677 (
            .O(N__28652),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv4 I__4676 (
            .O(N__28649),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__4675 (
            .O(N__28644),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__4674 (
            .O(N__28641),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__4673 (
            .O(N__28638),
            .I(N__28634));
    InMux I__4672 (
            .O(N__28637),
            .I(N__28631));
    LocalMux I__4671 (
            .O(N__28634),
            .I(N__28626));
    LocalMux I__4670 (
            .O(N__28631),
            .I(N__28626));
    Odrv12 I__4669 (
            .O(N__28626),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    CEMux I__4668 (
            .O(N__28623),
            .I(N__28605));
    CEMux I__4667 (
            .O(N__28622),
            .I(N__28605));
    CEMux I__4666 (
            .O(N__28621),
            .I(N__28605));
    CEMux I__4665 (
            .O(N__28620),
            .I(N__28605));
    CEMux I__4664 (
            .O(N__28619),
            .I(N__28605));
    CEMux I__4663 (
            .O(N__28618),
            .I(N__28605));
    GlobalMux I__4662 (
            .O(N__28605),
            .I(N__28602));
    gio2CtrlBuf I__4661 (
            .O(N__28602),
            .I(\delay_measurement_inst.delay_hc_timer.N_393_i_g ));
    InMux I__4660 (
            .O(N__28599),
            .I(N__28593));
    InMux I__4659 (
            .O(N__28598),
            .I(N__28593));
    LocalMux I__4658 (
            .O(N__28593),
            .I(N__28590));
    Odrv4 I__4657 (
            .O(N__28590),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__4656 (
            .O(N__28587),
            .I(N__28583));
    CascadeMux I__4655 (
            .O(N__28586),
            .I(N__28580));
    InMux I__4654 (
            .O(N__28583),
            .I(N__28575));
    InMux I__4653 (
            .O(N__28580),
            .I(N__28575));
    LocalMux I__4652 (
            .O(N__28575),
            .I(N__28572));
    Span4Mux_v I__4651 (
            .O(N__28572),
            .I(N__28568));
    InMux I__4650 (
            .O(N__28571),
            .I(N__28565));
    Span4Mux_h I__4649 (
            .O(N__28568),
            .I(N__28562));
    LocalMux I__4648 (
            .O(N__28565),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__4647 (
            .O(N__28562),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__4646 (
            .O(N__28557),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__4645 (
            .O(N__28554),
            .I(N__28551));
    InMux I__4644 (
            .O(N__28551),
            .I(N__28547));
    InMux I__4643 (
            .O(N__28550),
            .I(N__28544));
    LocalMux I__4642 (
            .O(N__28547),
            .I(N__28541));
    LocalMux I__4641 (
            .O(N__28544),
            .I(N__28538));
    Span4Mux_h I__4640 (
            .O(N__28541),
            .I(N__28532));
    Span4Mux_h I__4639 (
            .O(N__28538),
            .I(N__28532));
    InMux I__4638 (
            .O(N__28537),
            .I(N__28529));
    Span4Mux_v I__4637 (
            .O(N__28532),
            .I(N__28526));
    LocalMux I__4636 (
            .O(N__28529),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__4635 (
            .O(N__28526),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__4634 (
            .O(N__28521),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__4633 (
            .O(N__28518),
            .I(N__28515));
    InMux I__4632 (
            .O(N__28515),
            .I(N__28511));
    InMux I__4631 (
            .O(N__28514),
            .I(N__28508));
    LocalMux I__4630 (
            .O(N__28511),
            .I(N__28502));
    LocalMux I__4629 (
            .O(N__28508),
            .I(N__28502));
    InMux I__4628 (
            .O(N__28507),
            .I(N__28499));
    Span4Mux_v I__4627 (
            .O(N__28502),
            .I(N__28496));
    LocalMux I__4626 (
            .O(N__28499),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__4625 (
            .O(N__28496),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__4624 (
            .O(N__28491),
            .I(bfn_10_21_0_));
    InMux I__4623 (
            .O(N__28488),
            .I(N__28484));
    InMux I__4622 (
            .O(N__28487),
            .I(N__28481));
    LocalMux I__4621 (
            .O(N__28484),
            .I(N__28475));
    LocalMux I__4620 (
            .O(N__28481),
            .I(N__28475));
    InMux I__4619 (
            .O(N__28480),
            .I(N__28472));
    Span4Mux_v I__4618 (
            .O(N__28475),
            .I(N__28469));
    LocalMux I__4617 (
            .O(N__28472),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__4616 (
            .O(N__28469),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__4615 (
            .O(N__28464),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__4614 (
            .O(N__28461),
            .I(N__28454));
    InMux I__4613 (
            .O(N__28460),
            .I(N__28454));
    InMux I__4612 (
            .O(N__28459),
            .I(N__28451));
    LocalMux I__4611 (
            .O(N__28454),
            .I(N__28448));
    LocalMux I__4610 (
            .O(N__28451),
            .I(N__28443));
    Span4Mux_v I__4609 (
            .O(N__28448),
            .I(N__28443));
    Odrv4 I__4608 (
            .O(N__28443),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__4607 (
            .O(N__28440),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__4606 (
            .O(N__28437),
            .I(N__28433));
    CascadeMux I__4605 (
            .O(N__28436),
            .I(N__28430));
    InMux I__4604 (
            .O(N__28433),
            .I(N__28424));
    InMux I__4603 (
            .O(N__28430),
            .I(N__28424));
    InMux I__4602 (
            .O(N__28429),
            .I(N__28421));
    LocalMux I__4601 (
            .O(N__28424),
            .I(N__28418));
    LocalMux I__4600 (
            .O(N__28421),
            .I(N__28413));
    Span4Mux_v I__4599 (
            .O(N__28418),
            .I(N__28413));
    Odrv4 I__4598 (
            .O(N__28413),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__4597 (
            .O(N__28410),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__4596 (
            .O(N__28407),
            .I(N__28403));
    CascadeMux I__4595 (
            .O(N__28406),
            .I(N__28400));
    InMux I__4594 (
            .O(N__28403),
            .I(N__28395));
    InMux I__4593 (
            .O(N__28400),
            .I(N__28395));
    LocalMux I__4592 (
            .O(N__28395),
            .I(N__28391));
    InMux I__4591 (
            .O(N__28394),
            .I(N__28388));
    Span4Mux_v I__4590 (
            .O(N__28391),
            .I(N__28385));
    LocalMux I__4589 (
            .O(N__28388),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv4 I__4588 (
            .O(N__28385),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__4587 (
            .O(N__28380),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__4586 (
            .O(N__28377),
            .I(N__28374));
    InMux I__4585 (
            .O(N__28374),
            .I(N__28370));
    InMux I__4584 (
            .O(N__28373),
            .I(N__28367));
    LocalMux I__4583 (
            .O(N__28370),
            .I(N__28361));
    LocalMux I__4582 (
            .O(N__28367),
            .I(N__28361));
    InMux I__4581 (
            .O(N__28366),
            .I(N__28358));
    Span4Mux_v I__4580 (
            .O(N__28361),
            .I(N__28355));
    LocalMux I__4579 (
            .O(N__28358),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv4 I__4578 (
            .O(N__28355),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__4577 (
            .O(N__28350),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__4576 (
            .O(N__28347),
            .I(N__28344));
    InMux I__4575 (
            .O(N__28344),
            .I(N__28340));
    InMux I__4574 (
            .O(N__28343),
            .I(N__28337));
    LocalMux I__4573 (
            .O(N__28340),
            .I(N__28331));
    LocalMux I__4572 (
            .O(N__28337),
            .I(N__28331));
    InMux I__4571 (
            .O(N__28336),
            .I(N__28328));
    Span4Mux_v I__4570 (
            .O(N__28331),
            .I(N__28325));
    LocalMux I__4569 (
            .O(N__28328),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__4568 (
            .O(N__28325),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__4567 (
            .O(N__28320),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__4566 (
            .O(N__28317),
            .I(N__28311));
    InMux I__4565 (
            .O(N__28316),
            .I(N__28311));
    LocalMux I__4564 (
            .O(N__28311),
            .I(N__28307));
    InMux I__4563 (
            .O(N__28310),
            .I(N__28304));
    Span4Mux_v I__4562 (
            .O(N__28307),
            .I(N__28301));
    LocalMux I__4561 (
            .O(N__28304),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__4560 (
            .O(N__28301),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__4559 (
            .O(N__28296),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__4558 (
            .O(N__28293),
            .I(N__28286));
    InMux I__4557 (
            .O(N__28292),
            .I(N__28286));
    InMux I__4556 (
            .O(N__28291),
            .I(N__28283));
    LocalMux I__4555 (
            .O(N__28286),
            .I(N__28280));
    LocalMux I__4554 (
            .O(N__28283),
            .I(N__28275));
    Span4Mux_v I__4553 (
            .O(N__28280),
            .I(N__28275));
    Odrv4 I__4552 (
            .O(N__28275),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__4551 (
            .O(N__28272),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__4550 (
            .O(N__28269),
            .I(N__28265));
    CascadeMux I__4549 (
            .O(N__28268),
            .I(N__28262));
    InMux I__4548 (
            .O(N__28265),
            .I(N__28259));
    InMux I__4547 (
            .O(N__28262),
            .I(N__28256));
    LocalMux I__4546 (
            .O(N__28259),
            .I(N__28250));
    LocalMux I__4545 (
            .O(N__28256),
            .I(N__28250));
    InMux I__4544 (
            .O(N__28255),
            .I(N__28247));
    Span4Mux_v I__4543 (
            .O(N__28250),
            .I(N__28244));
    LocalMux I__4542 (
            .O(N__28247),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__4541 (
            .O(N__28244),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__4540 (
            .O(N__28239),
            .I(bfn_10_20_0_));
    CascadeMux I__4539 (
            .O(N__28236),
            .I(N__28233));
    InMux I__4538 (
            .O(N__28233),
            .I(N__28229));
    CascadeMux I__4537 (
            .O(N__28232),
            .I(N__28226));
    LocalMux I__4536 (
            .O(N__28229),
            .I(N__28222));
    InMux I__4535 (
            .O(N__28226),
            .I(N__28219));
    InMux I__4534 (
            .O(N__28225),
            .I(N__28216));
    Span4Mux_h I__4533 (
            .O(N__28222),
            .I(N__28211));
    LocalMux I__4532 (
            .O(N__28219),
            .I(N__28211));
    LocalMux I__4531 (
            .O(N__28216),
            .I(N__28206));
    Span4Mux_v I__4530 (
            .O(N__28211),
            .I(N__28206));
    Odrv4 I__4529 (
            .O(N__28206),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__4528 (
            .O(N__28203),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__4527 (
            .O(N__28200),
            .I(N__28197));
    InMux I__4526 (
            .O(N__28197),
            .I(N__28193));
    InMux I__4525 (
            .O(N__28196),
            .I(N__28190));
    LocalMux I__4524 (
            .O(N__28193),
            .I(N__28186));
    LocalMux I__4523 (
            .O(N__28190),
            .I(N__28183));
    InMux I__4522 (
            .O(N__28189),
            .I(N__28180));
    Span4Mux_h I__4521 (
            .O(N__28186),
            .I(N__28175));
    Span4Mux_h I__4520 (
            .O(N__28183),
            .I(N__28175));
    LocalMux I__4519 (
            .O(N__28180),
            .I(N__28170));
    Span4Mux_v I__4518 (
            .O(N__28175),
            .I(N__28170));
    Odrv4 I__4517 (
            .O(N__28170),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__4516 (
            .O(N__28167),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__4515 (
            .O(N__28164),
            .I(N__28158));
    InMux I__4514 (
            .O(N__28163),
            .I(N__28158));
    LocalMux I__4513 (
            .O(N__28158),
            .I(N__28155));
    Span4Mux_h I__4512 (
            .O(N__28155),
            .I(N__28151));
    InMux I__4511 (
            .O(N__28154),
            .I(N__28148));
    Span4Mux_v I__4510 (
            .O(N__28151),
            .I(N__28145));
    LocalMux I__4509 (
            .O(N__28148),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__4508 (
            .O(N__28145),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__4507 (
            .O(N__28140),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__4506 (
            .O(N__28137),
            .I(N__28131));
    InMux I__4505 (
            .O(N__28136),
            .I(N__28131));
    LocalMux I__4504 (
            .O(N__28131),
            .I(N__28127));
    InMux I__4503 (
            .O(N__28130),
            .I(N__28124));
    Span4Mux_v I__4502 (
            .O(N__28127),
            .I(N__28121));
    LocalMux I__4501 (
            .O(N__28124),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__4500 (
            .O(N__28121),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__4499 (
            .O(N__28116),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__4498 (
            .O(N__28113),
            .I(N__28109));
    CascadeMux I__4497 (
            .O(N__28112),
            .I(N__28106));
    InMux I__4496 (
            .O(N__28109),
            .I(N__28101));
    InMux I__4495 (
            .O(N__28106),
            .I(N__28101));
    LocalMux I__4494 (
            .O(N__28101),
            .I(N__28097));
    InMux I__4493 (
            .O(N__28100),
            .I(N__28094));
    Span4Mux_v I__4492 (
            .O(N__28097),
            .I(N__28091));
    LocalMux I__4491 (
            .O(N__28094),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__4490 (
            .O(N__28091),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__4489 (
            .O(N__28086),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__4488 (
            .O(N__28083),
            .I(N__28079));
    InMux I__4487 (
            .O(N__28082),
            .I(N__28074));
    LocalMux I__4486 (
            .O(N__28079),
            .I(N__28071));
    InMux I__4485 (
            .O(N__28078),
            .I(N__28068));
    InMux I__4484 (
            .O(N__28077),
            .I(N__28065));
    LocalMux I__4483 (
            .O(N__28074),
            .I(elapsed_time_ns_1_RNIMHKEE1_0_5));
    Odrv4 I__4482 (
            .O(N__28071),
            .I(elapsed_time_ns_1_RNIMHKEE1_0_5));
    LocalMux I__4481 (
            .O(N__28068),
            .I(elapsed_time_ns_1_RNIMHKEE1_0_5));
    LocalMux I__4480 (
            .O(N__28065),
            .I(elapsed_time_ns_1_RNIMHKEE1_0_5));
    CascadeMux I__4479 (
            .O(N__28056),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31_cascade_));
    InMux I__4478 (
            .O(N__28053),
            .I(N__28050));
    LocalMux I__4477 (
            .O(N__28050),
            .I(N__28046));
    InMux I__4476 (
            .O(N__28049),
            .I(N__28043));
    Span4Mux_h I__4475 (
            .O(N__28046),
            .I(N__28037));
    LocalMux I__4474 (
            .O(N__28043),
            .I(N__28037));
    InMux I__4473 (
            .O(N__28042),
            .I(N__28034));
    Span4Mux_v I__4472 (
            .O(N__28037),
            .I(N__28031));
    LocalMux I__4471 (
            .O(N__28034),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv4 I__4470 (
            .O(N__28031),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__4469 (
            .O(N__28026),
            .I(N__28022));
    InMux I__4468 (
            .O(N__28025),
            .I(N__28019));
    LocalMux I__4467 (
            .O(N__28022),
            .I(N__28016));
    LocalMux I__4466 (
            .O(N__28019),
            .I(N__28013));
    Span4Mux_v I__4465 (
            .O(N__28016),
            .I(N__28008));
    Span4Mux_v I__4464 (
            .O(N__28013),
            .I(N__28008));
    Odrv4 I__4463 (
            .O(N__28008),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__4462 (
            .O(N__28005),
            .I(N__28002));
    LocalMux I__4461 (
            .O(N__28002),
            .I(N__27998));
    InMux I__4460 (
            .O(N__28001),
            .I(N__27995));
    Span4Mux_v I__4459 (
            .O(N__27998),
            .I(N__27990));
    LocalMux I__4458 (
            .O(N__27995),
            .I(N__27990));
    Span4Mux_v I__4457 (
            .O(N__27990),
            .I(N__27986));
    InMux I__4456 (
            .O(N__27989),
            .I(N__27983));
    Odrv4 I__4455 (
            .O(N__27986),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__4454 (
            .O(N__27983),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    CascadeMux I__4453 (
            .O(N__27978),
            .I(N__27974));
    InMux I__4452 (
            .O(N__27977),
            .I(N__27971));
    InMux I__4451 (
            .O(N__27974),
            .I(N__27968));
    LocalMux I__4450 (
            .O(N__27971),
            .I(N__27965));
    LocalMux I__4449 (
            .O(N__27968),
            .I(N__27962));
    Span4Mux_v I__4448 (
            .O(N__27965),
            .I(N__27959));
    Span4Mux_v I__4447 (
            .O(N__27962),
            .I(N__27956));
    Odrv4 I__4446 (
            .O(N__27959),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__4445 (
            .O(N__27956),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__4444 (
            .O(N__27951),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__4443 (
            .O(N__27948),
            .I(N__27944));
    InMux I__4442 (
            .O(N__27947),
            .I(N__27941));
    InMux I__4441 (
            .O(N__27944),
            .I(N__27938));
    LocalMux I__4440 (
            .O(N__27941),
            .I(N__27932));
    LocalMux I__4439 (
            .O(N__27938),
            .I(N__27932));
    InMux I__4438 (
            .O(N__27937),
            .I(N__27929));
    Span4Mux_h I__4437 (
            .O(N__27932),
            .I(N__27926));
    LocalMux I__4436 (
            .O(N__27929),
            .I(N__27921));
    Span4Mux_v I__4435 (
            .O(N__27926),
            .I(N__27921));
    Odrv4 I__4434 (
            .O(N__27921),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    CascadeMux I__4433 (
            .O(N__27918),
            .I(N__27914));
    InMux I__4432 (
            .O(N__27917),
            .I(N__27911));
    InMux I__4431 (
            .O(N__27914),
            .I(N__27908));
    LocalMux I__4430 (
            .O(N__27911),
            .I(N__27905));
    LocalMux I__4429 (
            .O(N__27908),
            .I(N__27900));
    Span4Mux_h I__4428 (
            .O(N__27905),
            .I(N__27900));
    Odrv4 I__4427 (
            .O(N__27900),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__4426 (
            .O(N__27897),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__4425 (
            .O(N__27894),
            .I(N__27890));
    CascadeMux I__4424 (
            .O(N__27893),
            .I(N__27887));
    InMux I__4423 (
            .O(N__27890),
            .I(N__27882));
    InMux I__4422 (
            .O(N__27887),
            .I(N__27882));
    LocalMux I__4421 (
            .O(N__27882),
            .I(N__27879));
    Span4Mux_h I__4420 (
            .O(N__27879),
            .I(N__27875));
    InMux I__4419 (
            .O(N__27878),
            .I(N__27872));
    Span4Mux_v I__4418 (
            .O(N__27875),
            .I(N__27869));
    LocalMux I__4417 (
            .O(N__27872),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__4416 (
            .O(N__27869),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    CascadeMux I__4415 (
            .O(N__27864),
            .I(N__27861));
    InMux I__4414 (
            .O(N__27861),
            .I(N__27857));
    InMux I__4413 (
            .O(N__27860),
            .I(N__27854));
    LocalMux I__4412 (
            .O(N__27857),
            .I(N__27849));
    LocalMux I__4411 (
            .O(N__27854),
            .I(N__27849));
    Span4Mux_v I__4410 (
            .O(N__27849),
            .I(N__27846));
    Odrv4 I__4409 (
            .O(N__27846),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__4408 (
            .O(N__27843),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__4407 (
            .O(N__27840),
            .I(N__27836));
    CascadeMux I__4406 (
            .O(N__27839),
            .I(N__27833));
    InMux I__4405 (
            .O(N__27836),
            .I(N__27828));
    InMux I__4404 (
            .O(N__27833),
            .I(N__27828));
    LocalMux I__4403 (
            .O(N__27828),
            .I(N__27825));
    Span4Mux_h I__4402 (
            .O(N__27825),
            .I(N__27821));
    InMux I__4401 (
            .O(N__27824),
            .I(N__27818));
    Span4Mux_v I__4400 (
            .O(N__27821),
            .I(N__27815));
    LocalMux I__4399 (
            .O(N__27818),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__4398 (
            .O(N__27815),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__4397 (
            .O(N__27810),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__4396 (
            .O(N__27807),
            .I(N__27803));
    InMux I__4395 (
            .O(N__27806),
            .I(N__27800));
    LocalMux I__4394 (
            .O(N__27803),
            .I(elapsed_time_ns_1_RNI7JU8E1_0_24));
    LocalMux I__4393 (
            .O(N__27800),
            .I(elapsed_time_ns_1_RNI7JU8E1_0_24));
    InMux I__4392 (
            .O(N__27795),
            .I(N__27791));
    InMux I__4391 (
            .O(N__27794),
            .I(N__27788));
    LocalMux I__4390 (
            .O(N__27791),
            .I(elapsed_time_ns_1_RNIBNU8E1_0_28));
    LocalMux I__4389 (
            .O(N__27788),
            .I(elapsed_time_ns_1_RNIBNU8E1_0_28));
    CascadeMux I__4388 (
            .O(N__27783),
            .I(\delay_measurement_inst.delay_hc_timer.N_365_clk_cascade_ ));
    InMux I__4387 (
            .O(N__27780),
            .I(N__27773));
    InMux I__4386 (
            .O(N__27779),
            .I(N__27773));
    InMux I__4385 (
            .O(N__27778),
            .I(N__27770));
    LocalMux I__4384 (
            .O(N__27773),
            .I(\delay_measurement_inst.delay_hc_timer.N_367 ));
    LocalMux I__4383 (
            .O(N__27770),
            .I(\delay_measurement_inst.delay_hc_timer.N_367 ));
    CascadeMux I__4382 (
            .O(N__27765),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_ ));
    CascadeMux I__4381 (
            .O(N__27762),
            .I(N__27759));
    InMux I__4380 (
            .O(N__27759),
            .I(N__27755));
    InMux I__4379 (
            .O(N__27758),
            .I(N__27751));
    LocalMux I__4378 (
            .O(N__27755),
            .I(N__27748));
    InMux I__4377 (
            .O(N__27754),
            .I(N__27745));
    LocalMux I__4376 (
            .O(N__27751),
            .I(N__27735));
    Span4Mux_v I__4375 (
            .O(N__27748),
            .I(N__27735));
    LocalMux I__4374 (
            .O(N__27745),
            .I(N__27735));
    InMux I__4373 (
            .O(N__27744),
            .I(N__27731));
    InMux I__4372 (
            .O(N__27743),
            .I(N__27728));
    InMux I__4371 (
            .O(N__27742),
            .I(N__27725));
    Span4Mux_v I__4370 (
            .O(N__27735),
            .I(N__27722));
    InMux I__4369 (
            .O(N__27734),
            .I(N__27719));
    LocalMux I__4368 (
            .O(N__27731),
            .I(N__27714));
    LocalMux I__4367 (
            .O(N__27728),
            .I(N__27714));
    LocalMux I__4366 (
            .O(N__27725),
            .I(elapsed_time_ns_1_RNIDDC6P1_0_14));
    Odrv4 I__4365 (
            .O(N__27722),
            .I(elapsed_time_ns_1_RNIDDC6P1_0_14));
    LocalMux I__4364 (
            .O(N__27719),
            .I(elapsed_time_ns_1_RNIDDC6P1_0_14));
    Odrv4 I__4363 (
            .O(N__27714),
            .I(elapsed_time_ns_1_RNIDDC6P1_0_14));
    InMux I__4362 (
            .O(N__27705),
            .I(N__27702));
    LocalMux I__4361 (
            .O(N__27702),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14 ));
    CascadeMux I__4360 (
            .O(N__27699),
            .I(elapsed_time_ns_1_RNI6IU8E1_0_23_cascade_));
    CascadeMux I__4359 (
            .O(N__27696),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15_cascade_ ));
    InMux I__4358 (
            .O(N__27693),
            .I(N__27690));
    LocalMux I__4357 (
            .O(N__27690),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15 ));
    InMux I__4356 (
            .O(N__27687),
            .I(N__27684));
    LocalMux I__4355 (
            .O(N__27684),
            .I(N__27681));
    Odrv4 I__4354 (
            .O(N__27681),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1 ));
    CascadeMux I__4353 (
            .O(N__27678),
            .I(N__27675));
    InMux I__4352 (
            .O(N__27675),
            .I(N__27671));
    InMux I__4351 (
            .O(N__27674),
            .I(N__27668));
    LocalMux I__4350 (
            .O(N__27671),
            .I(elapsed_time_ns_1_RNI9LU8E1_0_26));
    LocalMux I__4349 (
            .O(N__27668),
            .I(elapsed_time_ns_1_RNI9LU8E1_0_26));
    CascadeMux I__4348 (
            .O(N__27663),
            .I(N__27660));
    InMux I__4347 (
            .O(N__27660),
            .I(N__27657));
    LocalMux I__4346 (
            .O(N__27657),
            .I(N__27654));
    Odrv12 I__4345 (
            .O(N__27654),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14 ));
    InMux I__4344 (
            .O(N__27651),
            .I(N__27648));
    LocalMux I__4343 (
            .O(N__27648),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20 ));
    CascadeMux I__4342 (
            .O(N__27645),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_ ));
    InMux I__4341 (
            .O(N__27642),
            .I(N__27638));
    InMux I__4340 (
            .O(N__27641),
            .I(N__27635));
    LocalMux I__4339 (
            .O(N__27638),
            .I(elapsed_time_ns_1_RNI5HU8E1_0_22));
    LocalMux I__4338 (
            .O(N__27635),
            .I(elapsed_time_ns_1_RNI5HU8E1_0_22));
    InMux I__4337 (
            .O(N__27630),
            .I(N__27622));
    InMux I__4336 (
            .O(N__27629),
            .I(N__27622));
    InMux I__4335 (
            .O(N__27628),
            .I(N__27619));
    InMux I__4334 (
            .O(N__27627),
            .I(N__27616));
    LocalMux I__4333 (
            .O(N__27622),
            .I(N__27613));
    LocalMux I__4332 (
            .O(N__27619),
            .I(N__27608));
    LocalMux I__4331 (
            .O(N__27616),
            .I(N__27608));
    Odrv4 I__4330 (
            .O(N__27613),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    Odrv4 I__4329 (
            .O(N__27608),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    CascadeMux I__4328 (
            .O(N__27603),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_ ));
    CascadeMux I__4327 (
            .O(N__27600),
            .I(\phase_controller_inst1.stoper_hc.N_326_cascade_ ));
    CascadeMux I__4326 (
            .O(N__27597),
            .I(N__27594));
    InMux I__4325 (
            .O(N__27594),
            .I(N__27591));
    LocalMux I__4324 (
            .O(N__27591),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ));
    CascadeMux I__4323 (
            .O(N__27588),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_ ));
    InMux I__4322 (
            .O(N__27585),
            .I(N__27582));
    LocalMux I__4321 (
            .O(N__27582),
            .I(N__27578));
    InMux I__4320 (
            .O(N__27581),
            .I(N__27575));
    Odrv4 I__4319 (
            .O(N__27578),
            .I(\phase_controller_inst1.stoper_hc.N_308 ));
    LocalMux I__4318 (
            .O(N__27575),
            .I(\phase_controller_inst1.stoper_hc.N_308 ));
    InMux I__4317 (
            .O(N__27570),
            .I(N__27566));
    InMux I__4316 (
            .O(N__27569),
            .I(N__27562));
    LocalMux I__4315 (
            .O(N__27566),
            .I(N__27559));
    CascadeMux I__4314 (
            .O(N__27565),
            .I(N__27556));
    LocalMux I__4313 (
            .O(N__27562),
            .I(N__27553));
    Span4Mux_h I__4312 (
            .O(N__27559),
            .I(N__27550));
    InMux I__4311 (
            .O(N__27556),
            .I(N__27547));
    Odrv4 I__4310 (
            .O(N__27553),
            .I(elapsed_time_ns_1_RNILGKEE1_0_4));
    Odrv4 I__4309 (
            .O(N__27550),
            .I(elapsed_time_ns_1_RNILGKEE1_0_4));
    LocalMux I__4308 (
            .O(N__27547),
            .I(elapsed_time_ns_1_RNILGKEE1_0_4));
    InMux I__4307 (
            .O(N__27540),
            .I(N__27537));
    LocalMux I__4306 (
            .O(N__27537),
            .I(elapsed_time_ns_1_RNIAMU8E1_0_27));
    CascadeMux I__4305 (
            .O(N__27534),
            .I(elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_));
    InMux I__4304 (
            .O(N__27531),
            .I(N__27528));
    LocalMux I__4303 (
            .O(N__27528),
            .I(elapsed_time_ns_1_RNI6IU8E1_0_23));
    CascadeMux I__4302 (
            .O(N__27525),
            .I(N__27509));
    CascadeMux I__4301 (
            .O(N__27524),
            .I(N__27506));
    CascadeMux I__4300 (
            .O(N__27523),
            .I(N__27503));
    InMux I__4299 (
            .O(N__27522),
            .I(N__27481));
    InMux I__4298 (
            .O(N__27521),
            .I(N__27481));
    InMux I__4297 (
            .O(N__27520),
            .I(N__27481));
    InMux I__4296 (
            .O(N__27519),
            .I(N__27481));
    InMux I__4295 (
            .O(N__27518),
            .I(N__27481));
    InMux I__4294 (
            .O(N__27517),
            .I(N__27481));
    InMux I__4293 (
            .O(N__27516),
            .I(N__27481));
    InMux I__4292 (
            .O(N__27515),
            .I(N__27478));
    InMux I__4291 (
            .O(N__27514),
            .I(N__27470));
    InMux I__4290 (
            .O(N__27513),
            .I(N__27459));
    InMux I__4289 (
            .O(N__27512),
            .I(N__27459));
    InMux I__4288 (
            .O(N__27509),
            .I(N__27459));
    InMux I__4287 (
            .O(N__27506),
            .I(N__27459));
    InMux I__4286 (
            .O(N__27503),
            .I(N__27459));
    InMux I__4285 (
            .O(N__27502),
            .I(N__27454));
    InMux I__4284 (
            .O(N__27501),
            .I(N__27454));
    InMux I__4283 (
            .O(N__27500),
            .I(N__27443));
    InMux I__4282 (
            .O(N__27499),
            .I(N__27443));
    InMux I__4281 (
            .O(N__27498),
            .I(N__27443));
    InMux I__4280 (
            .O(N__27497),
            .I(N__27443));
    InMux I__4279 (
            .O(N__27496),
            .I(N__27443));
    LocalMux I__4278 (
            .O(N__27481),
            .I(N__27440));
    LocalMux I__4277 (
            .O(N__27478),
            .I(N__27431));
    InMux I__4276 (
            .O(N__27477),
            .I(N__27420));
    InMux I__4275 (
            .O(N__27476),
            .I(N__27420));
    InMux I__4274 (
            .O(N__27475),
            .I(N__27420));
    InMux I__4273 (
            .O(N__27474),
            .I(N__27420));
    InMux I__4272 (
            .O(N__27473),
            .I(N__27420));
    LocalMux I__4271 (
            .O(N__27470),
            .I(N__27413));
    LocalMux I__4270 (
            .O(N__27459),
            .I(N__27413));
    LocalMux I__4269 (
            .O(N__27454),
            .I(N__27413));
    LocalMux I__4268 (
            .O(N__27443),
            .I(N__27408));
    Span4Mux_h I__4267 (
            .O(N__27440),
            .I(N__27408));
    InMux I__4266 (
            .O(N__27439),
            .I(N__27405));
    InMux I__4265 (
            .O(N__27438),
            .I(N__27394));
    InMux I__4264 (
            .O(N__27437),
            .I(N__27394));
    InMux I__4263 (
            .O(N__27436),
            .I(N__27394));
    InMux I__4262 (
            .O(N__27435),
            .I(N__27394));
    InMux I__4261 (
            .O(N__27434),
            .I(N__27394));
    Span4Mux_h I__4260 (
            .O(N__27431),
            .I(N__27391));
    LocalMux I__4259 (
            .O(N__27420),
            .I(N__27386));
    Span4Mux_v I__4258 (
            .O(N__27413),
            .I(N__27386));
    Span4Mux_v I__4257 (
            .O(N__27408),
            .I(N__27383));
    LocalMux I__4256 (
            .O(N__27405),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    LocalMux I__4255 (
            .O(N__27394),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__4254 (
            .O(N__27391),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__4253 (
            .O(N__27386),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__4252 (
            .O(N__27383),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    InMux I__4251 (
            .O(N__27372),
            .I(N__27362));
    InMux I__4250 (
            .O(N__27371),
            .I(N__27362));
    InMux I__4249 (
            .O(N__27370),
            .I(N__27362));
    InMux I__4248 (
            .O(N__27369),
            .I(N__27340));
    LocalMux I__4247 (
            .O(N__27362),
            .I(N__27337));
    InMux I__4246 (
            .O(N__27361),
            .I(N__27328));
    InMux I__4245 (
            .O(N__27360),
            .I(N__27328));
    InMux I__4244 (
            .O(N__27359),
            .I(N__27328));
    InMux I__4243 (
            .O(N__27358),
            .I(N__27328));
    CascadeMux I__4242 (
            .O(N__27357),
            .I(N__27325));
    InMux I__4241 (
            .O(N__27356),
            .I(N__27322));
    InMux I__4240 (
            .O(N__27355),
            .I(N__27319));
    InMux I__4239 (
            .O(N__27354),
            .I(N__27296));
    InMux I__4238 (
            .O(N__27353),
            .I(N__27296));
    InMux I__4237 (
            .O(N__27352),
            .I(N__27296));
    InMux I__4236 (
            .O(N__27351),
            .I(N__27296));
    InMux I__4235 (
            .O(N__27350),
            .I(N__27296));
    InMux I__4234 (
            .O(N__27349),
            .I(N__27296));
    InMux I__4233 (
            .O(N__27348),
            .I(N__27296));
    InMux I__4232 (
            .O(N__27347),
            .I(N__27285));
    InMux I__4231 (
            .O(N__27346),
            .I(N__27285));
    InMux I__4230 (
            .O(N__27345),
            .I(N__27285));
    InMux I__4229 (
            .O(N__27344),
            .I(N__27285));
    InMux I__4228 (
            .O(N__27343),
            .I(N__27285));
    LocalMux I__4227 (
            .O(N__27340),
            .I(N__27278));
    Span4Mux_v I__4226 (
            .O(N__27337),
            .I(N__27278));
    LocalMux I__4225 (
            .O(N__27328),
            .I(N__27278));
    InMux I__4224 (
            .O(N__27325),
            .I(N__27274));
    LocalMux I__4223 (
            .O(N__27322),
            .I(N__27271));
    LocalMux I__4222 (
            .O(N__27319),
            .I(N__27268));
    InMux I__4221 (
            .O(N__27318),
            .I(N__27263));
    InMux I__4220 (
            .O(N__27317),
            .I(N__27263));
    InMux I__4219 (
            .O(N__27316),
            .I(N__27260));
    InMux I__4218 (
            .O(N__27315),
            .I(N__27249));
    InMux I__4217 (
            .O(N__27314),
            .I(N__27249));
    InMux I__4216 (
            .O(N__27313),
            .I(N__27249));
    InMux I__4215 (
            .O(N__27312),
            .I(N__27249));
    InMux I__4214 (
            .O(N__27311),
            .I(N__27249));
    LocalMux I__4213 (
            .O(N__27296),
            .I(N__27244));
    LocalMux I__4212 (
            .O(N__27285),
            .I(N__27244));
    Span4Mux_v I__4211 (
            .O(N__27278),
            .I(N__27241));
    InMux I__4210 (
            .O(N__27277),
            .I(N__27238));
    LocalMux I__4209 (
            .O(N__27274),
            .I(N__27233));
    Span12Mux_s11_v I__4208 (
            .O(N__27271),
            .I(N__27233));
    Sp12to4 I__4207 (
            .O(N__27268),
            .I(N__27226));
    LocalMux I__4206 (
            .O(N__27263),
            .I(N__27226));
    LocalMux I__4205 (
            .O(N__27260),
            .I(N__27226));
    LocalMux I__4204 (
            .O(N__27249),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4203 (
            .O(N__27244),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__4202 (
            .O(N__27241),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__4201 (
            .O(N__27238),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__4200 (
            .O(N__27233),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__4199 (
            .O(N__27226),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    CascadeMux I__4198 (
            .O(N__27213),
            .I(N__27210));
    InMux I__4197 (
            .O(N__27210),
            .I(N__27207));
    LocalMux I__4196 (
            .O(N__27207),
            .I(N__27204));
    Span4Mux_v I__4195 (
            .O(N__27204),
            .I(N__27201));
    Odrv4 I__4194 (
            .O(N__27201),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__4193 (
            .O(N__27198),
            .I(N__27192));
    CascadeMux I__4192 (
            .O(N__27197),
            .I(N__27184));
    CascadeMux I__4191 (
            .O(N__27196),
            .I(N__27181));
    CascadeMux I__4190 (
            .O(N__27195),
            .I(N__27178));
    InMux I__4189 (
            .O(N__27192),
            .I(N__27171));
    CascadeMux I__4188 (
            .O(N__27191),
            .I(N__27157));
    CascadeMux I__4187 (
            .O(N__27190),
            .I(N__27154));
    CascadeMux I__4186 (
            .O(N__27189),
            .I(N__27151));
    InMux I__4185 (
            .O(N__27188),
            .I(N__27140));
    InMux I__4184 (
            .O(N__27187),
            .I(N__27140));
    InMux I__4183 (
            .O(N__27184),
            .I(N__27140));
    InMux I__4182 (
            .O(N__27181),
            .I(N__27140));
    InMux I__4181 (
            .O(N__27178),
            .I(N__27140));
    CascadeMux I__4180 (
            .O(N__27177),
            .I(N__27134));
    CascadeMux I__4179 (
            .O(N__27176),
            .I(N__27129));
    CascadeMux I__4178 (
            .O(N__27175),
            .I(N__27123));
    CascadeMux I__4177 (
            .O(N__27174),
            .I(N__27120));
    LocalMux I__4176 (
            .O(N__27171),
            .I(N__27117));
    InMux I__4175 (
            .O(N__27170),
            .I(N__27114));
    InMux I__4174 (
            .O(N__27169),
            .I(N__27111));
    InMux I__4173 (
            .O(N__27168),
            .I(N__27100));
    InMux I__4172 (
            .O(N__27167),
            .I(N__27100));
    InMux I__4171 (
            .O(N__27166),
            .I(N__27100));
    InMux I__4170 (
            .O(N__27165),
            .I(N__27100));
    InMux I__4169 (
            .O(N__27164),
            .I(N__27100));
    InMux I__4168 (
            .O(N__27163),
            .I(N__27085));
    InMux I__4167 (
            .O(N__27162),
            .I(N__27085));
    InMux I__4166 (
            .O(N__27161),
            .I(N__27085));
    InMux I__4165 (
            .O(N__27160),
            .I(N__27085));
    InMux I__4164 (
            .O(N__27157),
            .I(N__27085));
    InMux I__4163 (
            .O(N__27154),
            .I(N__27085));
    InMux I__4162 (
            .O(N__27151),
            .I(N__27085));
    LocalMux I__4161 (
            .O(N__27140),
            .I(N__27082));
    InMux I__4160 (
            .O(N__27139),
            .I(N__27071));
    InMux I__4159 (
            .O(N__27138),
            .I(N__27071));
    InMux I__4158 (
            .O(N__27137),
            .I(N__27071));
    InMux I__4157 (
            .O(N__27134),
            .I(N__27071));
    InMux I__4156 (
            .O(N__27133),
            .I(N__27071));
    InMux I__4155 (
            .O(N__27132),
            .I(N__27066));
    InMux I__4154 (
            .O(N__27129),
            .I(N__27066));
    InMux I__4153 (
            .O(N__27128),
            .I(N__27055));
    InMux I__4152 (
            .O(N__27127),
            .I(N__27055));
    InMux I__4151 (
            .O(N__27126),
            .I(N__27055));
    InMux I__4150 (
            .O(N__27123),
            .I(N__27055));
    InMux I__4149 (
            .O(N__27120),
            .I(N__27055));
    Span4Mux_v I__4148 (
            .O(N__27117),
            .I(N__27050));
    LocalMux I__4147 (
            .O(N__27114),
            .I(N__27050));
    LocalMux I__4146 (
            .O(N__27111),
            .I(N__27043));
    LocalMux I__4145 (
            .O(N__27100),
            .I(N__27043));
    LocalMux I__4144 (
            .O(N__27085),
            .I(N__27043));
    Span4Mux_v I__4143 (
            .O(N__27082),
            .I(N__27040));
    LocalMux I__4142 (
            .O(N__27071),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    LocalMux I__4141 (
            .O(N__27066),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    LocalMux I__4140 (
            .O(N__27055),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__4139 (
            .O(N__27050),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv12 I__4138 (
            .O(N__27043),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__4137 (
            .O(N__27040),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    InMux I__4136 (
            .O(N__27027),
            .I(N__27023));
    InMux I__4135 (
            .O(N__27026),
            .I(N__27019));
    LocalMux I__4134 (
            .O(N__27023),
            .I(N__27016));
    InMux I__4133 (
            .O(N__27022),
            .I(N__27013));
    LocalMux I__4132 (
            .O(N__27019),
            .I(N__27010));
    Span4Mux_h I__4131 (
            .O(N__27016),
            .I(N__27005));
    LocalMux I__4130 (
            .O(N__27013),
            .I(N__27002));
    Span4Mux_h I__4129 (
            .O(N__27010),
            .I(N__26999));
    InMux I__4128 (
            .O(N__27009),
            .I(N__26994));
    InMux I__4127 (
            .O(N__27008),
            .I(N__26994));
    Span4Mux_h I__4126 (
            .O(N__27005),
            .I(N__26991));
    Span12Mux_s11_v I__4125 (
            .O(N__27002),
            .I(N__26988));
    Sp12to4 I__4124 (
            .O(N__26999),
            .I(N__26983));
    LocalMux I__4123 (
            .O(N__26994),
            .I(N__26983));
    Odrv4 I__4122 (
            .O(N__26991),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv12 I__4121 (
            .O(N__26988),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv12 I__4120 (
            .O(N__26983),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__4119 (
            .O(N__26976),
            .I(N__26973));
    LocalMux I__4118 (
            .O(N__26973),
            .I(N__26970));
    Span4Mux_h I__4117 (
            .O(N__26970),
            .I(N__26967));
    Odrv4 I__4116 (
            .O(N__26967),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2 ));
    CascadeMux I__4115 (
            .O(N__26964),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_ ));
    CascadeMux I__4114 (
            .O(N__26961),
            .I(elapsed_time_ns_1_RNIJEKEE1_0_2_cascade_));
    InMux I__4113 (
            .O(N__26958),
            .I(N__26955));
    LocalMux I__4112 (
            .O(N__26955),
            .I(\phase_controller_inst1.stoper_hc.N_284 ));
    CascadeMux I__4111 (
            .O(N__26952),
            .I(N__26949));
    InMux I__4110 (
            .O(N__26949),
            .I(N__26943));
    InMux I__4109 (
            .O(N__26948),
            .I(N__26943));
    LocalMux I__4108 (
            .O(N__26943),
            .I(elapsed_time_ns_1_RNIJEKEE1_0_2));
    InMux I__4107 (
            .O(N__26940),
            .I(N__26934));
    InMux I__4106 (
            .O(N__26939),
            .I(N__26934));
    LocalMux I__4105 (
            .O(N__26934),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__4104 (
            .O(N__26931),
            .I(N__26927));
    InMux I__4103 (
            .O(N__26930),
            .I(N__26924));
    LocalMux I__4102 (
            .O(N__26927),
            .I(N__26916));
    LocalMux I__4101 (
            .O(N__26924),
            .I(N__26916));
    InMux I__4100 (
            .O(N__26923),
            .I(N__26911));
    InMux I__4099 (
            .O(N__26922),
            .I(N__26911));
    InMux I__4098 (
            .O(N__26921),
            .I(N__26908));
    Span4Mux_v I__4097 (
            .O(N__26916),
            .I(N__26905));
    LocalMux I__4096 (
            .O(N__26911),
            .I(elapsed_time_ns_1_RNI1I3CP1_0_9));
    LocalMux I__4095 (
            .O(N__26908),
            .I(elapsed_time_ns_1_RNI1I3CP1_0_9));
    Odrv4 I__4094 (
            .O(N__26905),
            .I(elapsed_time_ns_1_RNI1I3CP1_0_9));
    InMux I__4093 (
            .O(N__26898),
            .I(N__26893));
    InMux I__4092 (
            .O(N__26897),
            .I(N__26886));
    InMux I__4091 (
            .O(N__26896),
            .I(N__26886));
    LocalMux I__4090 (
            .O(N__26893),
            .I(N__26883));
    InMux I__4089 (
            .O(N__26892),
            .I(N__26878));
    InMux I__4088 (
            .O(N__26891),
            .I(N__26878));
    LocalMux I__4087 (
            .O(N__26886),
            .I(N__26875));
    Span4Mux_h I__4086 (
            .O(N__26883),
            .I(N__26872));
    LocalMux I__4085 (
            .O(N__26878),
            .I(N__26869));
    Span4Mux_v I__4084 (
            .O(N__26875),
            .I(N__26866));
    Odrv4 I__4083 (
            .O(N__26872),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv12 I__4082 (
            .O(N__26869),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__4081 (
            .O(N__26866),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__4080 (
            .O(N__26859),
            .I(N__26856));
    LocalMux I__4079 (
            .O(N__26856),
            .I(N__26853));
    Odrv4 I__4078 (
            .O(N__26853),
            .I(\current_shift_inst.PI_CTRL.integrator_i_21 ));
    CascadeMux I__4077 (
            .O(N__26850),
            .I(N__26847));
    InMux I__4076 (
            .O(N__26847),
            .I(N__26842));
    InMux I__4075 (
            .O(N__26846),
            .I(N__26839));
    InMux I__4074 (
            .O(N__26845),
            .I(N__26836));
    LocalMux I__4073 (
            .O(N__26842),
            .I(N__26833));
    LocalMux I__4072 (
            .O(N__26839),
            .I(N__26828));
    LocalMux I__4071 (
            .O(N__26836),
            .I(N__26825));
    Span4Mux_v I__4070 (
            .O(N__26833),
            .I(N__26822));
    InMux I__4069 (
            .O(N__26832),
            .I(N__26817));
    InMux I__4068 (
            .O(N__26831),
            .I(N__26817));
    Span4Mux_v I__4067 (
            .O(N__26828),
            .I(N__26812));
    Span4Mux_v I__4066 (
            .O(N__26825),
            .I(N__26812));
    Odrv4 I__4065 (
            .O(N__26822),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__4064 (
            .O(N__26817),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__4063 (
            .O(N__26812),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__4062 (
            .O(N__26805),
            .I(N__26802));
    InMux I__4061 (
            .O(N__26802),
            .I(N__26799));
    LocalMux I__4060 (
            .O(N__26799),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0 ));
    CascadeMux I__4059 (
            .O(N__26796),
            .I(N__26793));
    InMux I__4058 (
            .O(N__26793),
            .I(N__26790));
    LocalMux I__4057 (
            .O(N__26790),
            .I(N__26787));
    Span4Mux_h I__4056 (
            .O(N__26787),
            .I(N__26784));
    Odrv4 I__4055 (
            .O(N__26784),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10 ));
    InMux I__4054 (
            .O(N__26781),
            .I(N__26778));
    LocalMux I__4053 (
            .O(N__26778),
            .I(N__26775));
    Span4Mux_h I__4052 (
            .O(N__26775),
            .I(N__26772));
    Odrv4 I__4051 (
            .O(N__26772),
            .I(\current_shift_inst.PI_CTRL.integrator_i_6 ));
    InMux I__4050 (
            .O(N__26769),
            .I(N__26766));
    LocalMux I__4049 (
            .O(N__26766),
            .I(N__26763));
    Odrv4 I__4048 (
            .O(N__26763),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__4047 (
            .O(N__26760),
            .I(N__26756));
    CascadeMux I__4046 (
            .O(N__26759),
            .I(N__26752));
    InMux I__4045 (
            .O(N__26756),
            .I(N__26749));
    CascadeMux I__4044 (
            .O(N__26755),
            .I(N__26746));
    InMux I__4043 (
            .O(N__26752),
            .I(N__26743));
    LocalMux I__4042 (
            .O(N__26749),
            .I(N__26740));
    InMux I__4041 (
            .O(N__26746),
            .I(N__26737));
    LocalMux I__4040 (
            .O(N__26743),
            .I(N__26734));
    Span4Mux_v I__4039 (
            .O(N__26740),
            .I(N__26729));
    LocalMux I__4038 (
            .O(N__26737),
            .I(N__26729));
    Span4Mux_v I__4037 (
            .O(N__26734),
            .I(N__26722));
    Span4Mux_h I__4036 (
            .O(N__26729),
            .I(N__26722));
    InMux I__4035 (
            .O(N__26728),
            .I(N__26717));
    InMux I__4034 (
            .O(N__26727),
            .I(N__26717));
    Odrv4 I__4033 (
            .O(N__26722),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__4032 (
            .O(N__26717),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__4031 (
            .O(N__26712),
            .I(N__26709));
    InMux I__4030 (
            .O(N__26709),
            .I(N__26706));
    LocalMux I__4029 (
            .O(N__26706),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__4028 (
            .O(N__26703),
            .I(N__26700));
    LocalMux I__4027 (
            .O(N__26700),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__4026 (
            .O(N__26697),
            .I(N__26694));
    LocalMux I__4025 (
            .O(N__26694),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__4024 (
            .O(N__26691),
            .I(N__26687));
    InMux I__4023 (
            .O(N__26690),
            .I(N__26684));
    InMux I__4022 (
            .O(N__26687),
            .I(N__26679));
    LocalMux I__4021 (
            .O(N__26684),
            .I(N__26676));
    InMux I__4020 (
            .O(N__26683),
            .I(N__26673));
    InMux I__4019 (
            .O(N__26682),
            .I(N__26670));
    LocalMux I__4018 (
            .O(N__26679),
            .I(N__26667));
    Span4Mux_h I__4017 (
            .O(N__26676),
            .I(N__26664));
    LocalMux I__4016 (
            .O(N__26673),
            .I(N__26659));
    LocalMux I__4015 (
            .O(N__26670),
            .I(N__26659));
    Span4Mux_h I__4014 (
            .O(N__26667),
            .I(N__26654));
    Span4Mux_v I__4013 (
            .O(N__26664),
            .I(N__26654));
    Odrv12 I__4012 (
            .O(N__26659),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__4011 (
            .O(N__26654),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__4010 (
            .O(N__26649),
            .I(N__26646));
    InMux I__4009 (
            .O(N__26646),
            .I(N__26643));
    LocalMux I__4008 (
            .O(N__26643),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0 ));
    CascadeMux I__4007 (
            .O(N__26640),
            .I(N__26637));
    InMux I__4006 (
            .O(N__26637),
            .I(N__26633));
    InMux I__4005 (
            .O(N__26636),
            .I(N__26630));
    LocalMux I__4004 (
            .O(N__26633),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_14 ));
    LocalMux I__4003 (
            .O(N__26630),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_14 ));
    CascadeMux I__4002 (
            .O(N__26625),
            .I(N__26622));
    InMux I__4001 (
            .O(N__26622),
            .I(N__26619));
    LocalMux I__4000 (
            .O(N__26619),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0 ));
    CascadeMux I__3999 (
            .O(N__26616),
            .I(N__26613));
    InMux I__3998 (
            .O(N__26613),
            .I(N__26610));
    LocalMux I__3997 (
            .O(N__26610),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0 ));
    CascadeMux I__3996 (
            .O(N__26607),
            .I(N__26604));
    InMux I__3995 (
            .O(N__26604),
            .I(N__26601));
    LocalMux I__3994 (
            .O(N__26601),
            .I(N__26598));
    Odrv4 I__3993 (
            .O(N__26598),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0 ));
    CascadeMux I__3992 (
            .O(N__26595),
            .I(N__26592));
    InMux I__3991 (
            .O(N__26592),
            .I(N__26589));
    LocalMux I__3990 (
            .O(N__26589),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0 ));
    CascadeMux I__3989 (
            .O(N__26586),
            .I(N__26583));
    InMux I__3988 (
            .O(N__26583),
            .I(N__26580));
    LocalMux I__3987 (
            .O(N__26580),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0 ));
    CascadeMux I__3986 (
            .O(N__26577),
            .I(N__26574));
    InMux I__3985 (
            .O(N__26574),
            .I(N__26571));
    LocalMux I__3984 (
            .O(N__26571),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0 ));
    InMux I__3983 (
            .O(N__26568),
            .I(N__26564));
    CascadeMux I__3982 (
            .O(N__26567),
            .I(N__26561));
    LocalMux I__3981 (
            .O(N__26564),
            .I(N__26558));
    InMux I__3980 (
            .O(N__26561),
            .I(N__26555));
    Span4Mux_v I__3979 (
            .O(N__26558),
            .I(N__26550));
    LocalMux I__3978 (
            .O(N__26555),
            .I(N__26547));
    InMux I__3977 (
            .O(N__26554),
            .I(N__26543));
    InMux I__3976 (
            .O(N__26553),
            .I(N__26540));
    Span4Mux_v I__3975 (
            .O(N__26550),
            .I(N__26535));
    Span4Mux_h I__3974 (
            .O(N__26547),
            .I(N__26535));
    InMux I__3973 (
            .O(N__26546),
            .I(N__26532));
    LocalMux I__3972 (
            .O(N__26543),
            .I(N__26527));
    LocalMux I__3971 (
            .O(N__26540),
            .I(N__26527));
    Odrv4 I__3970 (
            .O(N__26535),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__3969 (
            .O(N__26532),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv12 I__3968 (
            .O(N__26527),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__3967 (
            .O(N__26520),
            .I(N__26517));
    InMux I__3966 (
            .O(N__26517),
            .I(N__26514));
    LocalMux I__3965 (
            .O(N__26514),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0 ));
    InMux I__3964 (
            .O(N__26511),
            .I(N__26506));
    InMux I__3963 (
            .O(N__26510),
            .I(N__26503));
    InMux I__3962 (
            .O(N__26509),
            .I(N__26500));
    LocalMux I__3961 (
            .O(N__26506),
            .I(N__26496));
    LocalMux I__3960 (
            .O(N__26503),
            .I(N__26493));
    LocalMux I__3959 (
            .O(N__26500),
            .I(N__26489));
    InMux I__3958 (
            .O(N__26499),
            .I(N__26486));
    Span4Mux_h I__3957 (
            .O(N__26496),
            .I(N__26481));
    Span4Mux_h I__3956 (
            .O(N__26493),
            .I(N__26481));
    InMux I__3955 (
            .O(N__26492),
            .I(N__26478));
    Span4Mux_h I__3954 (
            .O(N__26489),
            .I(N__26473));
    LocalMux I__3953 (
            .O(N__26486),
            .I(N__26473));
    Odrv4 I__3952 (
            .O(N__26481),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__3951 (
            .O(N__26478),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__3950 (
            .O(N__26473),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__3949 (
            .O(N__26466),
            .I(N__26463));
    InMux I__3948 (
            .O(N__26463),
            .I(N__26460));
    LocalMux I__3947 (
            .O(N__26460),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8 ));
    CascadeMux I__3946 (
            .O(N__26457),
            .I(N__26454));
    InMux I__3945 (
            .O(N__26454),
            .I(N__26451));
    LocalMux I__3944 (
            .O(N__26451),
            .I(N__26448));
    Span4Mux_h I__3943 (
            .O(N__26448),
            .I(N__26445));
    Odrv4 I__3942 (
            .O(N__26445),
            .I(\current_shift_inst.PI_CTRL.integrator_i_30 ));
    CascadeMux I__3941 (
            .O(N__26442),
            .I(N__26439));
    InMux I__3940 (
            .O(N__26439),
            .I(N__26436));
    LocalMux I__3939 (
            .O(N__26436),
            .I(N__26433));
    Odrv4 I__3938 (
            .O(N__26433),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6 ));
    CascadeMux I__3937 (
            .O(N__26430),
            .I(N__26427));
    InMux I__3936 (
            .O(N__26427),
            .I(N__26424));
    LocalMux I__3935 (
            .O(N__26424),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0 ));
    InMux I__3934 (
            .O(N__26421),
            .I(N__26417));
    CascadeMux I__3933 (
            .O(N__26420),
            .I(N__26412));
    LocalMux I__3932 (
            .O(N__26417),
            .I(N__26408));
    InMux I__3931 (
            .O(N__26416),
            .I(N__26405));
    InMux I__3930 (
            .O(N__26415),
            .I(N__26402));
    InMux I__3929 (
            .O(N__26412),
            .I(N__26399));
    InMux I__3928 (
            .O(N__26411),
            .I(N__26396));
    Span4Mux_h I__3927 (
            .O(N__26408),
            .I(N__26391));
    LocalMux I__3926 (
            .O(N__26405),
            .I(N__26391));
    LocalMux I__3925 (
            .O(N__26402),
            .I(N__26388));
    LocalMux I__3924 (
            .O(N__26399),
            .I(N__26385));
    LocalMux I__3923 (
            .O(N__26396),
            .I(N__26380));
    Span4Mux_v I__3922 (
            .O(N__26391),
            .I(N__26380));
    Odrv4 I__3921 (
            .O(N__26388),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__3920 (
            .O(N__26385),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__3919 (
            .O(N__26380),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__3918 (
            .O(N__26373),
            .I(N__26370));
    InMux I__3917 (
            .O(N__26370),
            .I(N__26367));
    LocalMux I__3916 (
            .O(N__26367),
            .I(N__26364));
    Odrv4 I__3915 (
            .O(N__26364),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0 ));
    InMux I__3914 (
            .O(N__26361),
            .I(N__26358));
    LocalMux I__3913 (
            .O(N__26358),
            .I(N__26354));
    InMux I__3912 (
            .O(N__26357),
            .I(N__26351));
    Span4Mux_h I__3911 (
            .O(N__26354),
            .I(N__26344));
    LocalMux I__3910 (
            .O(N__26351),
            .I(N__26344));
    InMux I__3909 (
            .O(N__26350),
            .I(N__26339));
    InMux I__3908 (
            .O(N__26349),
            .I(N__26339));
    Span4Mux_h I__3907 (
            .O(N__26344),
            .I(N__26335));
    LocalMux I__3906 (
            .O(N__26339),
            .I(N__26332));
    InMux I__3905 (
            .O(N__26338),
            .I(N__26329));
    Odrv4 I__3904 (
            .O(N__26335),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv12 I__3903 (
            .O(N__26332),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__3902 (
            .O(N__26329),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__3901 (
            .O(N__26322),
            .I(N__26319));
    InMux I__3900 (
            .O(N__26319),
            .I(N__26316));
    LocalMux I__3899 (
            .O(N__26316),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0 ));
    CascadeMux I__3898 (
            .O(N__26313),
            .I(N__26310));
    InMux I__3897 (
            .O(N__26310),
            .I(N__26307));
    LocalMux I__3896 (
            .O(N__26307),
            .I(N__26304));
    Odrv4 I__3895 (
            .O(N__26304),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0 ));
    CascadeMux I__3894 (
            .O(N__26301),
            .I(N__26295));
    InMux I__3893 (
            .O(N__26300),
            .I(N__26292));
    InMux I__3892 (
            .O(N__26299),
            .I(N__26288));
    InMux I__3891 (
            .O(N__26298),
            .I(N__26285));
    InMux I__3890 (
            .O(N__26295),
            .I(N__26282));
    LocalMux I__3889 (
            .O(N__26292),
            .I(N__26279));
    InMux I__3888 (
            .O(N__26291),
            .I(N__26276));
    LocalMux I__3887 (
            .O(N__26288),
            .I(N__26273));
    LocalMux I__3886 (
            .O(N__26285),
            .I(N__26268));
    LocalMux I__3885 (
            .O(N__26282),
            .I(N__26268));
    Span4Mux_h I__3884 (
            .O(N__26279),
            .I(N__26265));
    LocalMux I__3883 (
            .O(N__26276),
            .I(N__26260));
    Span4Mux_h I__3882 (
            .O(N__26273),
            .I(N__26260));
    Odrv12 I__3881 (
            .O(N__26268),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__3880 (
            .O(N__26265),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__3879 (
            .O(N__26260),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    CascadeMux I__3878 (
            .O(N__26253),
            .I(N__26250));
    InMux I__3877 (
            .O(N__26250),
            .I(N__26247));
    LocalMux I__3876 (
            .O(N__26247),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13 ));
    InMux I__3875 (
            .O(N__26244),
            .I(N__26241));
    LocalMux I__3874 (
            .O(N__26241),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    CascadeMux I__3873 (
            .O(N__26238),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0_cascade_ ));
    CascadeMux I__3872 (
            .O(N__26235),
            .I(N__26232));
    InMux I__3871 (
            .O(N__26232),
            .I(N__26229));
    LocalMux I__3870 (
            .O(N__26229),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4 ));
    InMux I__3869 (
            .O(N__26226),
            .I(N__26223));
    LocalMux I__3868 (
            .O(N__26223),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ));
    InMux I__3867 (
            .O(N__26220),
            .I(N__26217));
    LocalMux I__3866 (
            .O(N__26217),
            .I(\current_shift_inst.PI_CTRL.integrator_i_1 ));
    CascadeMux I__3865 (
            .O(N__26214),
            .I(N__26211));
    InMux I__3864 (
            .O(N__26211),
            .I(N__26208));
    LocalMux I__3863 (
            .O(N__26208),
            .I(N__26205));
    Span4Mux_v I__3862 (
            .O(N__26205),
            .I(N__26202));
    Span4Mux_h I__3861 (
            .O(N__26202),
            .I(N__26197));
    InMux I__3860 (
            .O(N__26201),
            .I(N__26192));
    InMux I__3859 (
            .O(N__26200),
            .I(N__26192));
    Odrv4 I__3858 (
            .O(N__26197),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__3857 (
            .O(N__26192),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__3856 (
            .O(N__26187),
            .I(N__26184));
    LocalMux I__3855 (
            .O(N__26184),
            .I(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ));
    CascadeMux I__3854 (
            .O(N__26181),
            .I(N__26178));
    InMux I__3853 (
            .O(N__26178),
            .I(N__26175));
    LocalMux I__3852 (
            .O(N__26175),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0 ));
    CascadeMux I__3851 (
            .O(N__26172),
            .I(N__26169));
    InMux I__3850 (
            .O(N__26169),
            .I(N__26163));
    InMux I__3849 (
            .O(N__26168),
            .I(N__26160));
    InMux I__3848 (
            .O(N__26167),
            .I(N__26157));
    InMux I__3847 (
            .O(N__26166),
            .I(N__26154));
    LocalMux I__3846 (
            .O(N__26163),
            .I(N__26151));
    LocalMux I__3845 (
            .O(N__26160),
            .I(N__26146));
    LocalMux I__3844 (
            .O(N__26157),
            .I(N__26146));
    LocalMux I__3843 (
            .O(N__26154),
            .I(N__26143));
    Span4Mux_v I__3842 (
            .O(N__26151),
            .I(N__26139));
    Span12Mux_s10_v I__3841 (
            .O(N__26146),
            .I(N__26136));
    Span4Mux_h I__3840 (
            .O(N__26143),
            .I(N__26133));
    InMux I__3839 (
            .O(N__26142),
            .I(N__26130));
    Odrv4 I__3838 (
            .O(N__26139),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv12 I__3837 (
            .O(N__26136),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__3836 (
            .O(N__26133),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__3835 (
            .O(N__26130),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    CascadeMux I__3834 (
            .O(N__26121),
            .I(N__26118));
    InMux I__3833 (
            .O(N__26118),
            .I(N__26115));
    LocalMux I__3832 (
            .O(N__26115),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12 ));
    InMux I__3831 (
            .O(N__26112),
            .I(N__26109));
    LocalMux I__3830 (
            .O(N__26109),
            .I(\current_shift_inst.PI_CTRL.integrator_i_10 ));
    InMux I__3829 (
            .O(N__26106),
            .I(N__26102));
    InMux I__3828 (
            .O(N__26105),
            .I(N__26099));
    LocalMux I__3827 (
            .O(N__26102),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__3826 (
            .O(N__26099),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__3825 (
            .O(N__26094),
            .I(N__26090));
    InMux I__3824 (
            .O(N__26093),
            .I(N__26087));
    LocalMux I__3823 (
            .O(N__26090),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__3822 (
            .O(N__26087),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__3821 (
            .O(N__26082),
            .I(N__26079));
    LocalMux I__3820 (
            .O(N__26079),
            .I(N__26076));
    Odrv4 I__3819 (
            .O(N__26076),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df28 ));
    InMux I__3818 (
            .O(N__26073),
            .I(N__26070));
    LocalMux I__3817 (
            .O(N__26070),
            .I(N__26067));
    Span4Mux_v I__3816 (
            .O(N__26067),
            .I(N__26064));
    Odrv4 I__3815 (
            .O(N__26064),
            .I(\current_shift_inst.PI_CTRL.integrator_i_9 ));
    InMux I__3814 (
            .O(N__26061),
            .I(N__26058));
    LocalMux I__3813 (
            .O(N__26058),
            .I(N__26055));
    Odrv12 I__3812 (
            .O(N__26055),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__3811 (
            .O(N__26052),
            .I(N__26049));
    LocalMux I__3810 (
            .O(N__26049),
            .I(N__26046));
    Odrv4 I__3809 (
            .O(N__26046),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    CascadeMux I__3808 (
            .O(N__26043),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_ ));
    InMux I__3807 (
            .O(N__26040),
            .I(N__26037));
    LocalMux I__3806 (
            .O(N__26037),
            .I(N__26034));
    Odrv4 I__3805 (
            .O(N__26034),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ));
    CascadeMux I__3804 (
            .O(N__26031),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ));
    CascadeMux I__3803 (
            .O(N__26028),
            .I(N__26025));
    InMux I__3802 (
            .O(N__26025),
            .I(N__26021));
    InMux I__3801 (
            .O(N__26024),
            .I(N__26017));
    LocalMux I__3800 (
            .O(N__26021),
            .I(N__26014));
    InMux I__3799 (
            .O(N__26020),
            .I(N__26009));
    LocalMux I__3798 (
            .O(N__26017),
            .I(N__26006));
    Span4Mux_h I__3797 (
            .O(N__26014),
            .I(N__26003));
    InMux I__3796 (
            .O(N__26013),
            .I(N__25998));
    InMux I__3795 (
            .O(N__26012),
            .I(N__25998));
    LocalMux I__3794 (
            .O(N__26009),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__3793 (
            .O(N__26006),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__3792 (
            .O(N__26003),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__3791 (
            .O(N__25998),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__3790 (
            .O(N__25989),
            .I(N__25986));
    LocalMux I__3789 (
            .O(N__25986),
            .I(\current_shift_inst.PI_CTRL.N_71 ));
    IoInMux I__3788 (
            .O(N__25983),
            .I(N__25980));
    LocalMux I__3787 (
            .O(N__25980),
            .I(N__25977));
    Span4Mux_s3_v I__3786 (
            .O(N__25977),
            .I(N__25974));
    Span4Mux_h I__3785 (
            .O(N__25974),
            .I(N__25971));
    Sp12to4 I__3784 (
            .O(N__25971),
            .I(N__25968));
    Span12Mux_s11_v I__3783 (
            .O(N__25968),
            .I(N__25965));
    Span12Mux_v I__3782 (
            .O(N__25965),
            .I(N__25962));
    Odrv12 I__3781 (
            .O(N__25962),
            .I(\pll_inst.red_c_i ));
    InMux I__3780 (
            .O(N__25959),
            .I(N__25956));
    LocalMux I__3779 (
            .O(N__25956),
            .I(N__25953));
    Span4Mux_v I__3778 (
            .O(N__25953),
            .I(N__25950));
    Odrv4 I__3777 (
            .O(N__25950),
            .I(\current_shift_inst.PI_CTRL.integrator_i_20 ));
    InMux I__3776 (
            .O(N__25947),
            .I(N__25944));
    LocalMux I__3775 (
            .O(N__25944),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    InMux I__3774 (
            .O(N__25941),
            .I(N__25937));
    InMux I__3773 (
            .O(N__25940),
            .I(N__25934));
    LocalMux I__3772 (
            .O(N__25937),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__3771 (
            .O(N__25934),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__3770 (
            .O(N__25929),
            .I(N__25925));
    InMux I__3769 (
            .O(N__25928),
            .I(N__25922));
    LocalMux I__3768 (
            .O(N__25925),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__3767 (
            .O(N__25922),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__3766 (
            .O(N__25917),
            .I(N__25914));
    LocalMux I__3765 (
            .O(N__25914),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df24 ));
    CascadeMux I__3764 (
            .O(N__25911),
            .I(N__25908));
    InMux I__3763 (
            .O(N__25908),
            .I(N__25905));
    LocalMux I__3762 (
            .O(N__25905),
            .I(N__25902));
    Span4Mux_v I__3761 (
            .O(N__25902),
            .I(N__25899));
    Odrv4 I__3760 (
            .O(N__25899),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    InMux I__3759 (
            .O(N__25896),
            .I(N__25891));
    InMux I__3758 (
            .O(N__25895),
            .I(N__25886));
    InMux I__3757 (
            .O(N__25894),
            .I(N__25886));
    LocalMux I__3756 (
            .O(N__25891),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__3755 (
            .O(N__25886),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__3754 (
            .O(N__25881),
            .I(N__25877));
    InMux I__3753 (
            .O(N__25880),
            .I(N__25873));
    InMux I__3752 (
            .O(N__25877),
            .I(N__25868));
    InMux I__3751 (
            .O(N__25876),
            .I(N__25868));
    LocalMux I__3750 (
            .O(N__25873),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__3749 (
            .O(N__25868),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__3748 (
            .O(N__25863),
            .I(N__25860));
    InMux I__3747 (
            .O(N__25860),
            .I(N__25857));
    LocalMux I__3746 (
            .O(N__25857),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    InMux I__3745 (
            .O(N__25854),
            .I(N__25850));
    InMux I__3744 (
            .O(N__25853),
            .I(N__25847));
    LocalMux I__3743 (
            .O(N__25850),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    LocalMux I__3742 (
            .O(N__25847),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__3741 (
            .O(N__25842),
            .I(N__25838));
    InMux I__3740 (
            .O(N__25841),
            .I(N__25835));
    LocalMux I__3739 (
            .O(N__25838),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    LocalMux I__3738 (
            .O(N__25835),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__3737 (
            .O(N__25830),
            .I(N__25827));
    LocalMux I__3736 (
            .O(N__25827),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df20 ));
    InMux I__3735 (
            .O(N__25824),
            .I(N__25819));
    InMux I__3734 (
            .O(N__25823),
            .I(N__25814));
    InMux I__3733 (
            .O(N__25822),
            .I(N__25814));
    LocalMux I__3732 (
            .O(N__25819),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    LocalMux I__3731 (
            .O(N__25814),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__3730 (
            .O(N__25809),
            .I(N__25805));
    InMux I__3729 (
            .O(N__25808),
            .I(N__25800));
    InMux I__3728 (
            .O(N__25805),
            .I(N__25800));
    LocalMux I__3727 (
            .O(N__25800),
            .I(N__25797));
    Span4Mux_v I__3726 (
            .O(N__25797),
            .I(N__25794));
    Odrv4 I__3725 (
            .O(N__25794),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__3724 (
            .O(N__25791),
            .I(N__25786));
    InMux I__3723 (
            .O(N__25790),
            .I(N__25781));
    InMux I__3722 (
            .O(N__25789),
            .I(N__25781));
    LocalMux I__3721 (
            .O(N__25786),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__3720 (
            .O(N__25781),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__3719 (
            .O(N__25776),
            .I(N__25773));
    LocalMux I__3718 (
            .O(N__25773),
            .I(N__25770));
    Odrv12 I__3717 (
            .O(N__25770),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    InMux I__3716 (
            .O(N__25767),
            .I(N__25763));
    InMux I__3715 (
            .O(N__25766),
            .I(N__25760));
    LocalMux I__3714 (
            .O(N__25763),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    LocalMux I__3713 (
            .O(N__25760),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__3712 (
            .O(N__25755),
            .I(N__25751));
    InMux I__3711 (
            .O(N__25754),
            .I(N__25748));
    LocalMux I__3710 (
            .O(N__25751),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    LocalMux I__3709 (
            .O(N__25748),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__3708 (
            .O(N__25743),
            .I(N__25740));
    LocalMux I__3707 (
            .O(N__25740),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df22 ));
    InMux I__3706 (
            .O(N__25737),
            .I(N__25733));
    InMux I__3705 (
            .O(N__25736),
            .I(N__25730));
    LocalMux I__3704 (
            .O(N__25733),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__3703 (
            .O(N__25730),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__3702 (
            .O(N__25725),
            .I(N__25721));
    InMux I__3701 (
            .O(N__25724),
            .I(N__25718));
    LocalMux I__3700 (
            .O(N__25721),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__3699 (
            .O(N__25718),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__3698 (
            .O(N__25713),
            .I(N__25710));
    LocalMux I__3697 (
            .O(N__25710),
            .I(N__25707));
    Odrv4 I__3696 (
            .O(N__25707),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df26 ));
    InMux I__3695 (
            .O(N__25704),
            .I(N__25701));
    LocalMux I__3694 (
            .O(N__25701),
            .I(N__25698));
    Odrv4 I__3693 (
            .O(N__25698),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__3692 (
            .O(N__25695),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ));
    InMux I__3691 (
            .O(N__25692),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    InMux I__3690 (
            .O(N__25689),
            .I(N__25685));
    InMux I__3689 (
            .O(N__25688),
            .I(N__25682));
    LocalMux I__3688 (
            .O(N__25685),
            .I(N__25679));
    LocalMux I__3687 (
            .O(N__25682),
            .I(N__25676));
    Span4Mux_v I__3686 (
            .O(N__25679),
            .I(N__25671));
    Span4Mux_h I__3685 (
            .O(N__25676),
            .I(N__25671));
    Odrv4 I__3684 (
            .O(N__25671),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    CascadeMux I__3683 (
            .O(N__25668),
            .I(N__25665));
    InMux I__3682 (
            .O(N__25665),
            .I(N__25660));
    InMux I__3681 (
            .O(N__25664),
            .I(N__25656));
    InMux I__3680 (
            .O(N__25663),
            .I(N__25653));
    LocalMux I__3679 (
            .O(N__25660),
            .I(N__25650));
    InMux I__3678 (
            .O(N__25659),
            .I(N__25647));
    LocalMux I__3677 (
            .O(N__25656),
            .I(N__25644));
    LocalMux I__3676 (
            .O(N__25653),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__3675 (
            .O(N__25650),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    LocalMux I__3674 (
            .O(N__25647),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv12 I__3673 (
            .O(N__25644),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__3672 (
            .O(N__25635),
            .I(N__25632));
    InMux I__3671 (
            .O(N__25632),
            .I(N__25627));
    InMux I__3670 (
            .O(N__25631),
            .I(N__25624));
    InMux I__3669 (
            .O(N__25630),
            .I(N__25621));
    LocalMux I__3668 (
            .O(N__25627),
            .I(N__25618));
    LocalMux I__3667 (
            .O(N__25624),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__3666 (
            .O(N__25621),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv12 I__3665 (
            .O(N__25618),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__3664 (
            .O(N__25611),
            .I(N__25608));
    LocalMux I__3663 (
            .O(N__25608),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    InMux I__3662 (
            .O(N__25605),
            .I(N__25601));
    InMux I__3661 (
            .O(N__25604),
            .I(N__25598));
    LocalMux I__3660 (
            .O(N__25601),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__3659 (
            .O(N__25598),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__3658 (
            .O(N__25593),
            .I(N__25590));
    InMux I__3657 (
            .O(N__25590),
            .I(N__25587));
    LocalMux I__3656 (
            .O(N__25587),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__3655 (
            .O(N__25584),
            .I(N__25581));
    InMux I__3654 (
            .O(N__25581),
            .I(N__25578));
    LocalMux I__3653 (
            .O(N__25578),
            .I(N__25575));
    Odrv4 I__3652 (
            .O(N__25575),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__3651 (
            .O(N__25572),
            .I(N__25568));
    InMux I__3650 (
            .O(N__25571),
            .I(N__25565));
    LocalMux I__3649 (
            .O(N__25568),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__3648 (
            .O(N__25565),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__3647 (
            .O(N__25560),
            .I(N__25557));
    LocalMux I__3646 (
            .O(N__25557),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__3645 (
            .O(N__25554),
            .I(N__25551));
    InMux I__3644 (
            .O(N__25551),
            .I(N__25548));
    LocalMux I__3643 (
            .O(N__25548),
            .I(N__25545));
    Odrv4 I__3642 (
            .O(N__25545),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__3641 (
            .O(N__25542),
            .I(N__25538));
    InMux I__3640 (
            .O(N__25541),
            .I(N__25535));
    LocalMux I__3639 (
            .O(N__25538),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__3638 (
            .O(N__25535),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__3637 (
            .O(N__25530),
            .I(N__25527));
    LocalMux I__3636 (
            .O(N__25527),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__3635 (
            .O(N__25524),
            .I(N__25521));
    LocalMux I__3634 (
            .O(N__25521),
            .I(N__25518));
    Odrv4 I__3633 (
            .O(N__25518),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__3632 (
            .O(N__25515),
            .I(N__25511));
    InMux I__3631 (
            .O(N__25514),
            .I(N__25508));
    LocalMux I__3630 (
            .O(N__25511),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__3629 (
            .O(N__25508),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__3628 (
            .O(N__25503),
            .I(N__25500));
    InMux I__3627 (
            .O(N__25500),
            .I(N__25497));
    LocalMux I__3626 (
            .O(N__25497),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__3625 (
            .O(N__25494),
            .I(N__25491));
    LocalMux I__3624 (
            .O(N__25491),
            .I(N__25488));
    Odrv4 I__3623 (
            .O(N__25488),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__3622 (
            .O(N__25485),
            .I(N__25481));
    InMux I__3621 (
            .O(N__25484),
            .I(N__25478));
    LocalMux I__3620 (
            .O(N__25481),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__3619 (
            .O(N__25478),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__3618 (
            .O(N__25473),
            .I(N__25470));
    InMux I__3617 (
            .O(N__25470),
            .I(N__25467));
    LocalMux I__3616 (
            .O(N__25467),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__3615 (
            .O(N__25464),
            .I(N__25461));
    InMux I__3614 (
            .O(N__25461),
            .I(N__25458));
    LocalMux I__3613 (
            .O(N__25458),
            .I(N__25455));
    Odrv12 I__3612 (
            .O(N__25455),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__3611 (
            .O(N__25452),
            .I(N__25448));
    InMux I__3610 (
            .O(N__25451),
            .I(N__25445));
    LocalMux I__3609 (
            .O(N__25448),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__3608 (
            .O(N__25445),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__3607 (
            .O(N__25440),
            .I(N__25437));
    LocalMux I__3606 (
            .O(N__25437),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__3605 (
            .O(N__25434),
            .I(N__25431));
    LocalMux I__3604 (
            .O(N__25431),
            .I(N__25428));
    Odrv12 I__3603 (
            .O(N__25428),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__3602 (
            .O(N__25425),
            .I(N__25422));
    InMux I__3601 (
            .O(N__25422),
            .I(N__25418));
    InMux I__3600 (
            .O(N__25421),
            .I(N__25415));
    LocalMux I__3599 (
            .O(N__25418),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__3598 (
            .O(N__25415),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__3597 (
            .O(N__25410),
            .I(N__25407));
    InMux I__3596 (
            .O(N__25407),
            .I(N__25404));
    LocalMux I__3595 (
            .O(N__25404),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__3594 (
            .O(N__25401),
            .I(N__25398));
    LocalMux I__3593 (
            .O(N__25398),
            .I(N__25395));
    Span12Mux_s9_v I__3592 (
            .O(N__25395),
            .I(N__25392));
    Odrv12 I__3591 (
            .O(N__25392),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__3590 (
            .O(N__25389),
            .I(N__25385));
    InMux I__3589 (
            .O(N__25388),
            .I(N__25382));
    LocalMux I__3588 (
            .O(N__25385),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__3587 (
            .O(N__25382),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__3586 (
            .O(N__25377),
            .I(N__25374));
    InMux I__3585 (
            .O(N__25374),
            .I(N__25371));
    LocalMux I__3584 (
            .O(N__25371),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__3583 (
            .O(N__25368),
            .I(N__25364));
    InMux I__3582 (
            .O(N__25367),
            .I(N__25361));
    LocalMux I__3581 (
            .O(N__25364),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__3580 (
            .O(N__25361),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__3579 (
            .O(N__25356),
            .I(N__25353));
    LocalMux I__3578 (
            .O(N__25353),
            .I(N__25350));
    Odrv12 I__3577 (
            .O(N__25350),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__3576 (
            .O(N__25347),
            .I(N__25344));
    InMux I__3575 (
            .O(N__25344),
            .I(N__25341));
    LocalMux I__3574 (
            .O(N__25341),
            .I(N__25338));
    Odrv4 I__3573 (
            .O(N__25338),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__3572 (
            .O(N__25335),
            .I(N__25332));
    LocalMux I__3571 (
            .O(N__25332),
            .I(N__25329));
    Span4Mux_v I__3570 (
            .O(N__25329),
            .I(N__25326));
    Span4Mux_v I__3569 (
            .O(N__25326),
            .I(N__25323));
    Odrv4 I__3568 (
            .O(N__25323),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    InMux I__3567 (
            .O(N__25320),
            .I(N__25316));
    InMux I__3566 (
            .O(N__25319),
            .I(N__25313));
    LocalMux I__3565 (
            .O(N__25316),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__3564 (
            .O(N__25313),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__3563 (
            .O(N__25308),
            .I(N__25305));
    InMux I__3562 (
            .O(N__25305),
            .I(N__25302));
    LocalMux I__3561 (
            .O(N__25302),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__3560 (
            .O(N__25299),
            .I(N__25296));
    LocalMux I__3559 (
            .O(N__25296),
            .I(N__25293));
    Span4Mux_v I__3558 (
            .O(N__25293),
            .I(N__25290));
    Span4Mux_h I__3557 (
            .O(N__25290),
            .I(N__25287));
    Odrv4 I__3556 (
            .O(N__25287),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__3555 (
            .O(N__25284),
            .I(N__25280));
    InMux I__3554 (
            .O(N__25283),
            .I(N__25277));
    LocalMux I__3553 (
            .O(N__25280),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__3552 (
            .O(N__25277),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__3551 (
            .O(N__25272),
            .I(N__25269));
    InMux I__3550 (
            .O(N__25269),
            .I(N__25266));
    LocalMux I__3549 (
            .O(N__25266),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__3548 (
            .O(N__25263),
            .I(N__25259));
    InMux I__3547 (
            .O(N__25262),
            .I(N__25256));
    LocalMux I__3546 (
            .O(N__25259),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__3545 (
            .O(N__25256),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__3544 (
            .O(N__25251),
            .I(N__25248));
    InMux I__3543 (
            .O(N__25248),
            .I(N__25245));
    LocalMux I__3542 (
            .O(N__25245),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__3541 (
            .O(N__25242),
            .I(N__25239));
    LocalMux I__3540 (
            .O(N__25239),
            .I(N__25236));
    Odrv4 I__3539 (
            .O(N__25236),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__3538 (
            .O(N__25233),
            .I(N__25229));
    InMux I__3537 (
            .O(N__25232),
            .I(N__25226));
    LocalMux I__3536 (
            .O(N__25229),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__3535 (
            .O(N__25226),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__3534 (
            .O(N__25221),
            .I(N__25218));
    InMux I__3533 (
            .O(N__25218),
            .I(N__25215));
    LocalMux I__3532 (
            .O(N__25215),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    CascadeMux I__3531 (
            .O(N__25212),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9_cascade_ ));
    InMux I__3530 (
            .O(N__25209),
            .I(N__25206));
    LocalMux I__3529 (
            .O(N__25206),
            .I(\phase_controller_inst1.stoper_hc.N_267_iZ0Z_1 ));
    CascadeMux I__3528 (
            .O(N__25203),
            .I(N__25198));
    InMux I__3527 (
            .O(N__25202),
            .I(N__25195));
    InMux I__3526 (
            .O(N__25201),
            .I(N__25192));
    InMux I__3525 (
            .O(N__25198),
            .I(N__25189));
    LocalMux I__3524 (
            .O(N__25195),
            .I(N__25186));
    LocalMux I__3523 (
            .O(N__25192),
            .I(N__25183));
    LocalMux I__3522 (
            .O(N__25189),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__3521 (
            .O(N__25186),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__3520 (
            .O(N__25183),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__3519 (
            .O(N__25176),
            .I(N__25173));
    LocalMux I__3518 (
            .O(N__25173),
            .I(N__25170));
    Span4Mux_v I__3517 (
            .O(N__25170),
            .I(N__25167));
    Odrv4 I__3516 (
            .O(N__25167),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__3515 (
            .O(N__25164),
            .I(N__25161));
    InMux I__3514 (
            .O(N__25161),
            .I(N__25158));
    LocalMux I__3513 (
            .O(N__25158),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__3512 (
            .O(N__25155),
            .I(N__25151));
    InMux I__3511 (
            .O(N__25154),
            .I(N__25148));
    LocalMux I__3510 (
            .O(N__25151),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__3509 (
            .O(N__25148),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__3508 (
            .O(N__25143),
            .I(N__25140));
    InMux I__3507 (
            .O(N__25140),
            .I(N__25137));
    LocalMux I__3506 (
            .O(N__25137),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__3505 (
            .O(N__25134),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9_cascade_ ));
    CascadeMux I__3504 (
            .O(N__25131),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i_cascade_ ));
    CascadeMux I__3503 (
            .O(N__25128),
            .I(elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_));
    InMux I__3502 (
            .O(N__25125),
            .I(N__25122));
    LocalMux I__3501 (
            .O(N__25122),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18 ));
    InMux I__3500 (
            .O(N__25119),
            .I(N__25116));
    LocalMux I__3499 (
            .O(N__25116),
            .I(N__25113));
    Span4Mux_v I__3498 (
            .O(N__25113),
            .I(N__25110));
    Odrv4 I__3497 (
            .O(N__25110),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17 ));
    InMux I__3496 (
            .O(N__25107),
            .I(N__25101));
    CascadeMux I__3495 (
            .O(N__25106),
            .I(N__25098));
    InMux I__3494 (
            .O(N__25105),
            .I(N__25093));
    InMux I__3493 (
            .O(N__25104),
            .I(N__25093));
    LocalMux I__3492 (
            .O(N__25101),
            .I(N__25090));
    InMux I__3491 (
            .O(N__25098),
            .I(N__25087));
    LocalMux I__3490 (
            .O(N__25093),
            .I(N__25084));
    Odrv4 I__3489 (
            .O(N__25090),
            .I(elapsed_time_ns_1_RNIFFC6P1_0_16));
    LocalMux I__3488 (
            .O(N__25087),
            .I(elapsed_time_ns_1_RNIFFC6P1_0_16));
    Odrv12 I__3487 (
            .O(N__25084),
            .I(elapsed_time_ns_1_RNIFFC6P1_0_16));
    CascadeMux I__3486 (
            .O(N__25077),
            .I(\phase_controller_inst1.stoper_hc.N_267_iZ0Z_1_cascade_ ));
    CascadeMux I__3485 (
            .O(N__25074),
            .I(elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_));
    InMux I__3484 (
            .O(N__25071),
            .I(N__25065));
    InMux I__3483 (
            .O(N__25070),
            .I(N__25065));
    LocalMux I__3482 (
            .O(N__25065),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    InMux I__3481 (
            .O(N__25062),
            .I(N__25056));
    InMux I__3480 (
            .O(N__25061),
            .I(N__25056));
    LocalMux I__3479 (
            .O(N__25056),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__3478 (
            .O(N__25053),
            .I(elapsed_time_ns_1_RNILGKEE1_0_4_cascade_));
    CascadeMux I__3477 (
            .O(N__25050),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_ ));
    CascadeMux I__3476 (
            .O(N__25047),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_ ));
    CascadeMux I__3475 (
            .O(N__25044),
            .I(elapsed_time_ns_1_RNIUE3CP1_0_6_cascade_));
    CascadeMux I__3474 (
            .O(N__25041),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ));
    InMux I__3473 (
            .O(N__25038),
            .I(N__25035));
    LocalMux I__3472 (
            .O(N__25035),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__3471 (
            .O(N__25032),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ));
    CascadeMux I__3470 (
            .O(N__25029),
            .I(N__25026));
    InMux I__3469 (
            .O(N__25026),
            .I(N__25023));
    LocalMux I__3468 (
            .O(N__25023),
            .I(N__25020));
    Odrv4 I__3467 (
            .O(N__25020),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__3466 (
            .O(N__25017),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ));
    InMux I__3465 (
            .O(N__25014),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ));
    InMux I__3464 (
            .O(N__25011),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ));
    InMux I__3463 (
            .O(N__25008),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ));
    InMux I__3462 (
            .O(N__25005),
            .I(bfn_9_13_0_));
    CascadeMux I__3461 (
            .O(N__25002),
            .I(N__24999));
    InMux I__3460 (
            .O(N__24999),
            .I(N__24996));
    LocalMux I__3459 (
            .O(N__24996),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__3458 (
            .O(N__24993),
            .I(N__24990));
    LocalMux I__3457 (
            .O(N__24990),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3 ));
    InMux I__3456 (
            .O(N__24987),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ));
    InMux I__3455 (
            .O(N__24984),
            .I(N__24981));
    LocalMux I__3454 (
            .O(N__24981),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__3453 (
            .O(N__24978),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ));
    InMux I__3452 (
            .O(N__24975),
            .I(N__24972));
    LocalMux I__3451 (
            .O(N__24972),
            .I(N__24969));
    Odrv4 I__3450 (
            .O(N__24969),
            .I(\current_shift_inst.PI_CTRL.integrator_i_19 ));
    CascadeMux I__3449 (
            .O(N__24966),
            .I(N__24963));
    InMux I__3448 (
            .O(N__24963),
            .I(N__24960));
    LocalMux I__3447 (
            .O(N__24960),
            .I(N__24957));
    Odrv12 I__3446 (
            .O(N__24957),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__3445 (
            .O(N__24954),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ));
    CascadeMux I__3444 (
            .O(N__24951),
            .I(N__24948));
    InMux I__3443 (
            .O(N__24948),
            .I(N__24945));
    LocalMux I__3442 (
            .O(N__24945),
            .I(N__24942));
    Odrv4 I__3441 (
            .O(N__24942),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__3440 (
            .O(N__24939),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ));
    CascadeMux I__3439 (
            .O(N__24936),
            .I(N__24933));
    InMux I__3438 (
            .O(N__24933),
            .I(N__24930));
    LocalMux I__3437 (
            .O(N__24930),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__3436 (
            .O(N__24927),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ));
    InMux I__3435 (
            .O(N__24924),
            .I(N__24921));
    LocalMux I__3434 (
            .O(N__24921),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__3433 (
            .O(N__24918),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ));
    InMux I__3432 (
            .O(N__24915),
            .I(N__24912));
    LocalMux I__3431 (
            .O(N__24912),
            .I(N__24909));
    Span4Mux_v I__3430 (
            .O(N__24909),
            .I(N__24906));
    Span4Mux_v I__3429 (
            .O(N__24906),
            .I(N__24903));
    Odrv4 I__3428 (
            .O(N__24903),
            .I(\current_shift_inst.PI_CTRL.integrator_i_23 ));
    InMux I__3427 (
            .O(N__24900),
            .I(N__24897));
    LocalMux I__3426 (
            .O(N__24897),
            .I(N__24894));
    Odrv4 I__3425 (
            .O(N__24894),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__3424 (
            .O(N__24891),
            .I(bfn_9_12_0_));
    InMux I__3423 (
            .O(N__24888),
            .I(N__24885));
    LocalMux I__3422 (
            .O(N__24885),
            .I(N__24882));
    Odrv4 I__3421 (
            .O(N__24882),
            .I(\current_shift_inst.PI_CTRL.integrator_i_24 ));
    CascadeMux I__3420 (
            .O(N__24879),
            .I(N__24876));
    InMux I__3419 (
            .O(N__24876),
            .I(N__24873));
    LocalMux I__3418 (
            .O(N__24873),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__3417 (
            .O(N__24870),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ));
    CascadeMux I__3416 (
            .O(N__24867),
            .I(N__24864));
    InMux I__3415 (
            .O(N__24864),
            .I(N__24861));
    LocalMux I__3414 (
            .O(N__24861),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__3413 (
            .O(N__24858),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ));
    CascadeMux I__3412 (
            .O(N__24855),
            .I(N__24852));
    InMux I__3411 (
            .O(N__24852),
            .I(N__24849));
    LocalMux I__3410 (
            .O(N__24849),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__3409 (
            .O(N__24846),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ));
    InMux I__3408 (
            .O(N__24843),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ));
    CascadeMux I__3407 (
            .O(N__24840),
            .I(N__24837));
    InMux I__3406 (
            .O(N__24837),
            .I(N__24834));
    LocalMux I__3405 (
            .O(N__24834),
            .I(N__24831));
    Odrv4 I__3404 (
            .O(N__24831),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__3403 (
            .O(N__24828),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ));
    InMux I__3402 (
            .O(N__24825),
            .I(N__24822));
    LocalMux I__3401 (
            .O(N__24822),
            .I(N__24819));
    Odrv4 I__3400 (
            .O(N__24819),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__3399 (
            .O(N__24816),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ));
    CascadeMux I__3398 (
            .O(N__24813),
            .I(N__24810));
    InMux I__3397 (
            .O(N__24810),
            .I(N__24807));
    LocalMux I__3396 (
            .O(N__24807),
            .I(N__24804));
    Odrv4 I__3395 (
            .O(N__24804),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__3394 (
            .O(N__24801),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ));
    InMux I__3393 (
            .O(N__24798),
            .I(N__24795));
    LocalMux I__3392 (
            .O(N__24795),
            .I(N__24792));
    Odrv4 I__3391 (
            .O(N__24792),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__3390 (
            .O(N__24789),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ));
    InMux I__3389 (
            .O(N__24786),
            .I(N__24783));
    LocalMux I__3388 (
            .O(N__24783),
            .I(N__24780));
    Odrv12 I__3387 (
            .O(N__24780),
            .I(\current_shift_inst.PI_CTRL.integrator_i_15 ));
    CascadeMux I__3386 (
            .O(N__24777),
            .I(N__24774));
    InMux I__3385 (
            .O(N__24774),
            .I(N__24771));
    LocalMux I__3384 (
            .O(N__24771),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__3383 (
            .O(N__24768),
            .I(bfn_9_11_0_));
    InMux I__3382 (
            .O(N__24765),
            .I(N__24762));
    LocalMux I__3381 (
            .O(N__24762),
            .I(N__24759));
    Odrv4 I__3380 (
            .O(N__24759),
            .I(\current_shift_inst.PI_CTRL.integrator_i_16 ));
    CascadeMux I__3379 (
            .O(N__24756),
            .I(N__24753));
    InMux I__3378 (
            .O(N__24753),
            .I(N__24750));
    LocalMux I__3377 (
            .O(N__24750),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0 ));
    InMux I__3376 (
            .O(N__24747),
            .I(N__24744));
    LocalMux I__3375 (
            .O(N__24744),
            .I(N__24741));
    Span4Mux_v I__3374 (
            .O(N__24741),
            .I(N__24738));
    Odrv4 I__3373 (
            .O(N__24738),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__3372 (
            .O(N__24735),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ));
    CascadeMux I__3371 (
            .O(N__24732),
            .I(N__24729));
    InMux I__3370 (
            .O(N__24729),
            .I(N__24726));
    LocalMux I__3369 (
            .O(N__24726),
            .I(N__24723));
    Span4Mux_v I__3368 (
            .O(N__24723),
            .I(N__24720));
    Odrv4 I__3367 (
            .O(N__24720),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__3366 (
            .O(N__24717),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ));
    InMux I__3365 (
            .O(N__24714),
            .I(N__24711));
    LocalMux I__3364 (
            .O(N__24711),
            .I(N__24708));
    Odrv4 I__3363 (
            .O(N__24708),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__3362 (
            .O(N__24705),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ));
    InMux I__3361 (
            .O(N__24702),
            .I(N__24699));
    LocalMux I__3360 (
            .O(N__24699),
            .I(\current_shift_inst.PI_CTRL.integrator_i_3 ));
    CascadeMux I__3359 (
            .O(N__24696),
            .I(N__24693));
    InMux I__3358 (
            .O(N__24693),
            .I(N__24690));
    LocalMux I__3357 (
            .O(N__24690),
            .I(\current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7 ));
    InMux I__3356 (
            .O(N__24687),
            .I(N__24684));
    LocalMux I__3355 (
            .O(N__24684),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__3354 (
            .O(N__24681),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ));
    InMux I__3353 (
            .O(N__24678),
            .I(N__24675));
    LocalMux I__3352 (
            .O(N__24675),
            .I(N__24672));
    Odrv12 I__3351 (
            .O(N__24672),
            .I(\current_shift_inst.PI_CTRL.integrator_i_4 ));
    InMux I__3350 (
            .O(N__24669),
            .I(N__24666));
    LocalMux I__3349 (
            .O(N__24666),
            .I(N__24663));
    Odrv4 I__3348 (
            .O(N__24663),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__3347 (
            .O(N__24660),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ));
    InMux I__3346 (
            .O(N__24657),
            .I(N__24654));
    LocalMux I__3345 (
            .O(N__24654),
            .I(N__24651));
    Span4Mux_h I__3344 (
            .O(N__24651),
            .I(N__24648));
    Odrv4 I__3343 (
            .O(N__24648),
            .I(\current_shift_inst.PI_CTRL.integrator_i_5 ));
    CascadeMux I__3342 (
            .O(N__24645),
            .I(N__24642));
    InMux I__3341 (
            .O(N__24642),
            .I(N__24639));
    LocalMux I__3340 (
            .O(N__24639),
            .I(N__24636));
    Odrv4 I__3339 (
            .O(N__24636),
            .I(\current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9 ));
    InMux I__3338 (
            .O(N__24633),
            .I(N__24630));
    LocalMux I__3337 (
            .O(N__24630),
            .I(N__24627));
    Odrv4 I__3336 (
            .O(N__24627),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__3335 (
            .O(N__24624),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ));
    InMux I__3334 (
            .O(N__24621),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ));
    InMux I__3333 (
            .O(N__24618),
            .I(N__24615));
    LocalMux I__3332 (
            .O(N__24615),
            .I(\current_shift_inst.PI_CTRL.integrator_i_7 ));
    CascadeMux I__3331 (
            .O(N__24612),
            .I(N__24609));
    InMux I__3330 (
            .O(N__24609),
            .I(N__24606));
    LocalMux I__3329 (
            .O(N__24606),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11 ));
    InMux I__3328 (
            .O(N__24603),
            .I(N__24600));
    LocalMux I__3327 (
            .O(N__24600),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__3326 (
            .O(N__24597),
            .I(bfn_9_10_0_));
    InMux I__3325 (
            .O(N__24594),
            .I(N__24591));
    LocalMux I__3324 (
            .O(N__24591),
            .I(\current_shift_inst.PI_CTRL.integrator_i_8 ));
    InMux I__3323 (
            .O(N__24588),
            .I(N__24585));
    LocalMux I__3322 (
            .O(N__24585),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__3321 (
            .O(N__24582),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ));
    InMux I__3320 (
            .O(N__24579),
            .I(N__24576));
    LocalMux I__3319 (
            .O(N__24576),
            .I(N__24573));
    Odrv4 I__3318 (
            .O(N__24573),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ));
    InMux I__3317 (
            .O(N__24570),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ));
    InMux I__3316 (
            .O(N__24567),
            .I(N__24564));
    LocalMux I__3315 (
            .O(N__24564),
            .I(N__24561));
    Span4Mux_h I__3314 (
            .O(N__24561),
            .I(N__24555));
    InMux I__3313 (
            .O(N__24560),
            .I(N__24552));
    CascadeMux I__3312 (
            .O(N__24559),
            .I(N__24549));
    CascadeMux I__3311 (
            .O(N__24558),
            .I(N__24546));
    Sp12to4 I__3310 (
            .O(N__24555),
            .I(N__24543));
    LocalMux I__3309 (
            .O(N__24552),
            .I(N__24540));
    InMux I__3308 (
            .O(N__24549),
            .I(N__24535));
    InMux I__3307 (
            .O(N__24546),
            .I(N__24535));
    Span12Mux_s10_v I__3306 (
            .O(N__24543),
            .I(N__24532));
    Span4Mux_h I__3305 (
            .O(N__24540),
            .I(N__24529));
    LocalMux I__3304 (
            .O(N__24535),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__3303 (
            .O(N__24532),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__3302 (
            .O(N__24529),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    IoInMux I__3301 (
            .O(N__24522),
            .I(N__24519));
    LocalMux I__3300 (
            .O(N__24519),
            .I(s3_phy_c));
    InMux I__3299 (
            .O(N__24516),
            .I(N__24513));
    LocalMux I__3298 (
            .O(N__24513),
            .I(N__24510));
    Odrv12 I__3297 (
            .O(N__24510),
            .I(il_min_comp1_c));
    InMux I__3296 (
            .O(N__24507),
            .I(N__24504));
    LocalMux I__3295 (
            .O(N__24504),
            .I(N__24500));
    InMux I__3294 (
            .O(N__24503),
            .I(N__24497));
    Span4Mux_h I__3293 (
            .O(N__24500),
            .I(N__24490));
    LocalMux I__3292 (
            .O(N__24497),
            .I(N__24490));
    InMux I__3291 (
            .O(N__24496),
            .I(N__24487));
    InMux I__3290 (
            .O(N__24495),
            .I(N__24484));
    Span4Mux_v I__3289 (
            .O(N__24490),
            .I(N__24481));
    LocalMux I__3288 (
            .O(N__24487),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__3287 (
            .O(N__24484),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__3286 (
            .O(N__24481),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    ClkMux I__3285 (
            .O(N__24474),
            .I(N__24468));
    ClkMux I__3284 (
            .O(N__24473),
            .I(N__24468));
    GlobalMux I__3283 (
            .O(N__24468),
            .I(N__24465));
    gio2CtrlBuf I__3282 (
            .O(N__24465),
            .I(delay_hc_input_c_g));
    InMux I__3281 (
            .O(N__24462),
            .I(N__24459));
    LocalMux I__3280 (
            .O(N__24459),
            .I(N__24456));
    Span4Mux_v I__3279 (
            .O(N__24456),
            .I(N__24453));
    Span4Mux_h I__3278 (
            .O(N__24453),
            .I(N__24450));
    Odrv4 I__3277 (
            .O(N__24450),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__3276 (
            .O(N__24447),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__3275 (
            .O(N__24444),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__3274 (
            .O(N__24441),
            .I(bfn_8_26_0_));
    InMux I__3273 (
            .O(N__24438),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__3272 (
            .O(N__24435),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__3271 (
            .O(N__24432),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__3270 (
            .O(N__24429),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__3269 (
            .O(N__24426),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__3268 (
            .O(N__24423),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__3267 (
            .O(N__24420),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__3266 (
            .O(N__24417),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__3265 (
            .O(N__24414),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__3264 (
            .O(N__24411),
            .I(bfn_8_25_0_));
    InMux I__3263 (
            .O(N__24408),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__3262 (
            .O(N__24405),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__3261 (
            .O(N__24402),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__3260 (
            .O(N__24399),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__3259 (
            .O(N__24396),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__3258 (
            .O(N__24393),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__3257 (
            .O(N__24390),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__3256 (
            .O(N__24387),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__3255 (
            .O(N__24384),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__3254 (
            .O(N__24381),
            .I(bfn_8_24_0_));
    InMux I__3253 (
            .O(N__24378),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__3252 (
            .O(N__24375),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__3251 (
            .O(N__24372),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__3250 (
            .O(N__24369),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    CascadeMux I__3249 (
            .O(N__24366),
            .I(N__24363));
    InMux I__3248 (
            .O(N__24363),
            .I(N__24359));
    InMux I__3247 (
            .O(N__24362),
            .I(N__24356));
    LocalMux I__3246 (
            .O(N__24359),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__3245 (
            .O(N__24356),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    InMux I__3244 (
            .O(N__24351),
            .I(N__24347));
    InMux I__3243 (
            .O(N__24350),
            .I(N__24344));
    LocalMux I__3242 (
            .O(N__24347),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__3241 (
            .O(N__24344),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    InMux I__3240 (
            .O(N__24339),
            .I(N__24336));
    LocalMux I__3239 (
            .O(N__24336),
            .I(N__24329));
    InMux I__3238 (
            .O(N__24335),
            .I(N__24324));
    InMux I__3237 (
            .O(N__24334),
            .I(N__24324));
    InMux I__3236 (
            .O(N__24333),
            .I(N__24319));
    InMux I__3235 (
            .O(N__24332),
            .I(N__24319));
    Odrv4 I__3234 (
            .O(N__24329),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__3233 (
            .O(N__24324),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__3232 (
            .O(N__24319),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__3231 (
            .O(N__24312),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__3230 (
            .O(N__24309),
            .I(N__24306));
    InMux I__3229 (
            .O(N__24306),
            .I(N__24303));
    LocalMux I__3228 (
            .O(N__24303),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    InMux I__3227 (
            .O(N__24300),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__3226 (
            .O(N__24297),
            .I(N__24294));
    LocalMux I__3225 (
            .O(N__24294),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28 ));
    InMux I__3224 (
            .O(N__24291),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__3223 (
            .O(N__24288),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__3222 (
            .O(N__24285),
            .I(bfn_8_18_0_));
    InMux I__3221 (
            .O(N__24282),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__3220 (
            .O(N__24279),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__3219 (
            .O(N__24276),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__3218 (
            .O(N__24273),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__3217 (
            .O(N__24270),
            .I(N__24232));
    InMux I__3216 (
            .O(N__24269),
            .I(N__24232));
    InMux I__3215 (
            .O(N__24268),
            .I(N__24232));
    InMux I__3214 (
            .O(N__24267),
            .I(N__24232));
    InMux I__3213 (
            .O(N__24266),
            .I(N__24223));
    InMux I__3212 (
            .O(N__24265),
            .I(N__24223));
    InMux I__3211 (
            .O(N__24264),
            .I(N__24223));
    InMux I__3210 (
            .O(N__24263),
            .I(N__24223));
    InMux I__3209 (
            .O(N__24262),
            .I(N__24218));
    InMux I__3208 (
            .O(N__24261),
            .I(N__24218));
    InMux I__3207 (
            .O(N__24260),
            .I(N__24209));
    InMux I__3206 (
            .O(N__24259),
            .I(N__24209));
    InMux I__3205 (
            .O(N__24258),
            .I(N__24209));
    InMux I__3204 (
            .O(N__24257),
            .I(N__24209));
    InMux I__3203 (
            .O(N__24256),
            .I(N__24200));
    InMux I__3202 (
            .O(N__24255),
            .I(N__24200));
    InMux I__3201 (
            .O(N__24254),
            .I(N__24200));
    InMux I__3200 (
            .O(N__24253),
            .I(N__24200));
    InMux I__3199 (
            .O(N__24252),
            .I(N__24191));
    InMux I__3198 (
            .O(N__24251),
            .I(N__24191));
    InMux I__3197 (
            .O(N__24250),
            .I(N__24191));
    InMux I__3196 (
            .O(N__24249),
            .I(N__24191));
    InMux I__3195 (
            .O(N__24248),
            .I(N__24182));
    InMux I__3194 (
            .O(N__24247),
            .I(N__24182));
    InMux I__3193 (
            .O(N__24246),
            .I(N__24182));
    InMux I__3192 (
            .O(N__24245),
            .I(N__24182));
    InMux I__3191 (
            .O(N__24244),
            .I(N__24173));
    InMux I__3190 (
            .O(N__24243),
            .I(N__24173));
    InMux I__3189 (
            .O(N__24242),
            .I(N__24173));
    InMux I__3188 (
            .O(N__24241),
            .I(N__24173));
    LocalMux I__3187 (
            .O(N__24232),
            .I(N__24162));
    LocalMux I__3186 (
            .O(N__24223),
            .I(N__24162));
    LocalMux I__3185 (
            .O(N__24218),
            .I(N__24162));
    LocalMux I__3184 (
            .O(N__24209),
            .I(N__24162));
    LocalMux I__3183 (
            .O(N__24200),
            .I(N__24162));
    LocalMux I__3182 (
            .O(N__24191),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__3181 (
            .O(N__24182),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__3180 (
            .O(N__24173),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__3179 (
            .O(N__24162),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__3178 (
            .O(N__24153),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CEMux I__3177 (
            .O(N__24150),
            .I(N__24147));
    LocalMux I__3176 (
            .O(N__24147),
            .I(N__24141));
    CEMux I__3175 (
            .O(N__24146),
            .I(N__24138));
    CEMux I__3174 (
            .O(N__24145),
            .I(N__24135));
    CEMux I__3173 (
            .O(N__24144),
            .I(N__24132));
    Span4Mux_v I__3172 (
            .O(N__24141),
            .I(N__24129));
    LocalMux I__3171 (
            .O(N__24138),
            .I(N__24126));
    LocalMux I__3170 (
            .O(N__24135),
            .I(N__24123));
    LocalMux I__3169 (
            .O(N__24132),
            .I(N__24120));
    Span4Mux_h I__3168 (
            .O(N__24129),
            .I(N__24113));
    Span4Mux_v I__3167 (
            .O(N__24126),
            .I(N__24113));
    Span4Mux_h I__3166 (
            .O(N__24123),
            .I(N__24113));
    Odrv12 I__3165 (
            .O(N__24120),
            .I(\delay_measurement_inst.delay_hc_timer.N_394_i ));
    Odrv4 I__3164 (
            .O(N__24113),
            .I(\delay_measurement_inst.delay_hc_timer.N_394_i ));
    InMux I__3163 (
            .O(N__24108),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__3162 (
            .O(N__24105),
            .I(bfn_8_17_0_));
    InMux I__3161 (
            .O(N__24102),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__3160 (
            .O(N__24099),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__3159 (
            .O(N__24096),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__3158 (
            .O(N__24093),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__3157 (
            .O(N__24090),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__3156 (
            .O(N__24087),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__3155 (
            .O(N__24084),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__3154 (
            .O(N__24081),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__3153 (
            .O(N__24078),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__3152 (
            .O(N__24075),
            .I(bfn_8_16_0_));
    InMux I__3151 (
            .O(N__24072),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__3150 (
            .O(N__24069),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__3149 (
            .O(N__24066),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__3148 (
            .O(N__24063),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__3147 (
            .O(N__24060),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__3146 (
            .O(N__24057),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__3145 (
            .O(N__24054),
            .I(N__24046));
    InMux I__3144 (
            .O(N__24053),
            .I(N__24046));
    InMux I__3143 (
            .O(N__24052),
            .I(N__24043));
    InMux I__3142 (
            .O(N__24051),
            .I(N__24040));
    LocalMux I__3141 (
            .O(N__24046),
            .I(N__24037));
    LocalMux I__3140 (
            .O(N__24043),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__3139 (
            .O(N__24040),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__3138 (
            .O(N__24037),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__3137 (
            .O(N__24030),
            .I(N__24025));
    InMux I__3136 (
            .O(N__24029),
            .I(N__24022));
    InMux I__3135 (
            .O(N__24028),
            .I(N__24019));
    LocalMux I__3134 (
            .O(N__24025),
            .I(N__24016));
    LocalMux I__3133 (
            .O(N__24022),
            .I(N__24009));
    LocalMux I__3132 (
            .O(N__24019),
            .I(N__24009));
    Span4Mux_v I__3131 (
            .O(N__24016),
            .I(N__24009));
    Span4Mux_v I__3130 (
            .O(N__24009),
            .I(N__24006));
    Odrv4 I__3129 (
            .O(N__24006),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    CascadeMux I__3128 (
            .O(N__24003),
            .I(N__24000));
    InMux I__3127 (
            .O(N__24000),
            .I(N__23996));
    InMux I__3126 (
            .O(N__23999),
            .I(N__23993));
    LocalMux I__3125 (
            .O(N__23996),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__3124 (
            .O(N__23993),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__3123 (
            .O(N__23988),
            .I(N__23984));
    InMux I__3122 (
            .O(N__23987),
            .I(N__23981));
    LocalMux I__3121 (
            .O(N__23984),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    LocalMux I__3120 (
            .O(N__23981),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    InMux I__3119 (
            .O(N__23976),
            .I(bfn_8_15_0_));
    InMux I__3118 (
            .O(N__23973),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__3117 (
            .O(N__23970),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__3116 (
            .O(N__23967),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__3115 (
            .O(N__23964),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__3114 (
            .O(N__23961),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    CascadeMux I__3113 (
            .O(N__23958),
            .I(N__23955));
    InMux I__3112 (
            .O(N__23955),
            .I(N__23952));
    LocalMux I__3111 (
            .O(N__23952),
            .I(N__23949));
    Odrv12 I__3110 (
            .O(N__23949),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__3109 (
            .O(N__23946),
            .I(N__23943));
    InMux I__3108 (
            .O(N__23943),
            .I(N__23938));
    InMux I__3107 (
            .O(N__23942),
            .I(N__23935));
    InMux I__3106 (
            .O(N__23941),
            .I(N__23932));
    LocalMux I__3105 (
            .O(N__23938),
            .I(N__23928));
    LocalMux I__3104 (
            .O(N__23935),
            .I(N__23925));
    LocalMux I__3103 (
            .O(N__23932),
            .I(N__23922));
    InMux I__3102 (
            .O(N__23931),
            .I(N__23918));
    Span4Mux_v I__3101 (
            .O(N__23928),
            .I(N__23911));
    Span4Mux_v I__3100 (
            .O(N__23925),
            .I(N__23911));
    Span4Mux_v I__3099 (
            .O(N__23922),
            .I(N__23911));
    InMux I__3098 (
            .O(N__23921),
            .I(N__23908));
    LocalMux I__3097 (
            .O(N__23918),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__3096 (
            .O(N__23911),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__3095 (
            .O(N__23908),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    CascadeMux I__3094 (
            .O(N__23901),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20_cascade_ ));
    CascadeMux I__3093 (
            .O(N__23898),
            .I(N__23887));
    CascadeMux I__3092 (
            .O(N__23897),
            .I(N__23883));
    CascadeMux I__3091 (
            .O(N__23896),
            .I(N__23879));
    CascadeMux I__3090 (
            .O(N__23895),
            .I(N__23875));
    CascadeMux I__3089 (
            .O(N__23894),
            .I(N__23871));
    CascadeMux I__3088 (
            .O(N__23893),
            .I(N__23867));
    CascadeMux I__3087 (
            .O(N__23892),
            .I(N__23863));
    InMux I__3086 (
            .O(N__23891),
            .I(N__23844));
    InMux I__3085 (
            .O(N__23890),
            .I(N__23844));
    InMux I__3084 (
            .O(N__23887),
            .I(N__23844));
    InMux I__3083 (
            .O(N__23886),
            .I(N__23844));
    InMux I__3082 (
            .O(N__23883),
            .I(N__23844));
    InMux I__3081 (
            .O(N__23882),
            .I(N__23844));
    InMux I__3080 (
            .O(N__23879),
            .I(N__23844));
    InMux I__3079 (
            .O(N__23878),
            .I(N__23844));
    InMux I__3078 (
            .O(N__23875),
            .I(N__23827));
    InMux I__3077 (
            .O(N__23874),
            .I(N__23827));
    InMux I__3076 (
            .O(N__23871),
            .I(N__23827));
    InMux I__3075 (
            .O(N__23870),
            .I(N__23827));
    InMux I__3074 (
            .O(N__23867),
            .I(N__23827));
    InMux I__3073 (
            .O(N__23866),
            .I(N__23827));
    InMux I__3072 (
            .O(N__23863),
            .I(N__23827));
    InMux I__3071 (
            .O(N__23862),
            .I(N__23827));
    CascadeMux I__3070 (
            .O(N__23861),
            .I(N__23824));
    LocalMux I__3069 (
            .O(N__23844),
            .I(N__23818));
    LocalMux I__3068 (
            .O(N__23827),
            .I(N__23818));
    InMux I__3067 (
            .O(N__23824),
            .I(N__23813));
    InMux I__3066 (
            .O(N__23823),
            .I(N__23813));
    Span12Mux_v I__3065 (
            .O(N__23818),
            .I(N__23808));
    LocalMux I__3064 (
            .O(N__23813),
            .I(N__23808));
    Odrv12 I__3063 (
            .O(N__23808),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__3062 (
            .O(N__23805),
            .I(N__23802));
    InMux I__3061 (
            .O(N__23802),
            .I(N__23798));
    InMux I__3060 (
            .O(N__23801),
            .I(N__23794));
    LocalMux I__3059 (
            .O(N__23798),
            .I(N__23791));
    InMux I__3058 (
            .O(N__23797),
            .I(N__23788));
    LocalMux I__3057 (
            .O(N__23794),
            .I(N__23783));
    Span4Mux_v I__3056 (
            .O(N__23791),
            .I(N__23780));
    LocalMux I__3055 (
            .O(N__23788),
            .I(N__23777));
    InMux I__3054 (
            .O(N__23787),
            .I(N__23772));
    InMux I__3053 (
            .O(N__23786),
            .I(N__23772));
    Odrv4 I__3052 (
            .O(N__23783),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__3051 (
            .O(N__23780),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv12 I__3050 (
            .O(N__23777),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__3049 (
            .O(N__23772),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__3048 (
            .O(N__23763),
            .I(N__23760));
    LocalMux I__3047 (
            .O(N__23760),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__3046 (
            .O(N__23757),
            .I(N__23754));
    LocalMux I__3045 (
            .O(N__23754),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    CascadeMux I__3044 (
            .O(N__23751),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13_cascade_ ));
    CascadeMux I__3043 (
            .O(N__23748),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ));
    InMux I__3042 (
            .O(N__23745),
            .I(N__23742));
    LocalMux I__3041 (
            .O(N__23742),
            .I(\current_shift_inst.PI_CTRL.N_72 ));
    InMux I__3040 (
            .O(N__23739),
            .I(N__23736));
    LocalMux I__3039 (
            .O(N__23736),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    CascadeMux I__3038 (
            .O(N__23733),
            .I(N__23730));
    InMux I__3037 (
            .O(N__23730),
            .I(N__23726));
    InMux I__3036 (
            .O(N__23729),
            .I(N__23722));
    LocalMux I__3035 (
            .O(N__23726),
            .I(N__23717));
    InMux I__3034 (
            .O(N__23725),
            .I(N__23714));
    LocalMux I__3033 (
            .O(N__23722),
            .I(N__23711));
    InMux I__3032 (
            .O(N__23721),
            .I(N__23706));
    InMux I__3031 (
            .O(N__23720),
            .I(N__23706));
    Odrv12 I__3030 (
            .O(N__23717),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__3029 (
            .O(N__23714),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__3028 (
            .O(N__23711),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__3027 (
            .O(N__23706),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    CascadeMux I__3026 (
            .O(N__23697),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ));
    CascadeMux I__3025 (
            .O(N__23694),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12_cascade_ ));
    InMux I__3024 (
            .O(N__23691),
            .I(N__23688));
    LocalMux I__3023 (
            .O(N__23688),
            .I(N__23685));
    Odrv4 I__3022 (
            .O(N__23685),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ));
    InMux I__3021 (
            .O(N__23682),
            .I(N__23679));
    LocalMux I__3020 (
            .O(N__23679),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__3019 (
            .O(N__23676),
            .I(N__23673));
    LocalMux I__3018 (
            .O(N__23673),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ));
    InMux I__3017 (
            .O(N__23670),
            .I(N__23667));
    LocalMux I__3016 (
            .O(N__23667),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    InMux I__3015 (
            .O(N__23664),
            .I(N__23661));
    LocalMux I__3014 (
            .O(N__23661),
            .I(\phase_controller_inst2.start_timer_hc_RNO_0_0 ));
    InMux I__3013 (
            .O(N__23658),
            .I(N__23655));
    LocalMux I__3012 (
            .O(N__23655),
            .I(N__23652));
    Odrv4 I__3011 (
            .O(N__23652),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    CascadeMux I__3010 (
            .O(N__23649),
            .I(N__23646));
    InMux I__3009 (
            .O(N__23646),
            .I(N__23638));
    InMux I__3008 (
            .O(N__23645),
            .I(N__23638));
    InMux I__3007 (
            .O(N__23644),
            .I(N__23635));
    InMux I__3006 (
            .O(N__23643),
            .I(N__23632));
    LocalMux I__3005 (
            .O(N__23638),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__3004 (
            .O(N__23635),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__3003 (
            .O(N__23632),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__3002 (
            .O(N__23625),
            .I(N__23622));
    LocalMux I__3001 (
            .O(N__23622),
            .I(N__23618));
    InMux I__3000 (
            .O(N__23621),
            .I(N__23615));
    Span4Mux_s1_v I__2999 (
            .O(N__23618),
            .I(N__23610));
    LocalMux I__2998 (
            .O(N__23615),
            .I(N__23610));
    Span4Mux_v I__2997 (
            .O(N__23610),
            .I(N__23605));
    InMux I__2996 (
            .O(N__23609),
            .I(N__23602));
    InMux I__2995 (
            .O(N__23608),
            .I(N__23599));
    Span4Mux_h I__2994 (
            .O(N__23605),
            .I(N__23596));
    LocalMux I__2993 (
            .O(N__23602),
            .I(N__23591));
    LocalMux I__2992 (
            .O(N__23599),
            .I(N__23591));
    Sp12to4 I__2991 (
            .O(N__23596),
            .I(N__23588));
    Span4Mux_v I__2990 (
            .O(N__23591),
            .I(N__23585));
    Span12Mux_v I__2989 (
            .O(N__23588),
            .I(N__23582));
    Sp12to4 I__2988 (
            .O(N__23585),
            .I(N__23579));
    Span12Mux_v I__2987 (
            .O(N__23582),
            .I(N__23576));
    Span12Mux_h I__2986 (
            .O(N__23579),
            .I(N__23573));
    Span12Mux_h I__2985 (
            .O(N__23576),
            .I(N__23570));
    Span12Mux_v I__2984 (
            .O(N__23573),
            .I(N__23567));
    Odrv12 I__2983 (
            .O(N__23570),
            .I(start_stop_c));
    Odrv12 I__2982 (
            .O(N__23567),
            .I(start_stop_c));
    InMux I__2981 (
            .O(N__23562),
            .I(N__23559));
    LocalMux I__2980 (
            .O(N__23559),
            .I(N__23555));
    InMux I__2979 (
            .O(N__23558),
            .I(N__23550));
    Span12Mux_s6_v I__2978 (
            .O(N__23555),
            .I(N__23547));
    InMux I__2977 (
            .O(N__23554),
            .I(N__23542));
    InMux I__2976 (
            .O(N__23553),
            .I(N__23542));
    LocalMux I__2975 (
            .O(N__23550),
            .I(N__23539));
    Odrv12 I__2974 (
            .O(N__23547),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__2973 (
            .O(N__23542),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__2972 (
            .O(N__23539),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    IoInMux I__2971 (
            .O(N__23532),
            .I(N__23529));
    LocalMux I__2970 (
            .O(N__23529),
            .I(N__23526));
    Span4Mux_s3_v I__2969 (
            .O(N__23526),
            .I(N__23523));
    Odrv4 I__2968 (
            .O(N__23523),
            .I(s4_phy_c));
    InMux I__2967 (
            .O(N__23520),
            .I(N__23517));
    LocalMux I__2966 (
            .O(N__23517),
            .I(N__23514));
    Odrv12 I__2965 (
            .O(N__23514),
            .I(il_max_comp1_c));
    InMux I__2964 (
            .O(N__23511),
            .I(N__23508));
    LocalMux I__2963 (
            .O(N__23508),
            .I(il_max_comp1_D1));
    InMux I__2962 (
            .O(N__23505),
            .I(N__23498));
    InMux I__2961 (
            .O(N__23504),
            .I(N__23498));
    InMux I__2960 (
            .O(N__23503),
            .I(N__23495));
    LocalMux I__2959 (
            .O(N__23498),
            .I(N__23492));
    LocalMux I__2958 (
            .O(N__23495),
            .I(N__23489));
    Odrv4 I__2957 (
            .O(N__23492),
            .I(il_max_comp2_D2));
    Odrv4 I__2956 (
            .O(N__23489),
            .I(il_max_comp2_D2));
    InMux I__2955 (
            .O(N__23484),
            .I(N__23478));
    InMux I__2954 (
            .O(N__23483),
            .I(N__23478));
    LocalMux I__2953 (
            .O(N__23478),
            .I(N__23474));
    InMux I__2952 (
            .O(N__23477),
            .I(N__23471));
    Odrv4 I__2951 (
            .O(N__23474),
            .I(il_min_comp2_D2));
    LocalMux I__2950 (
            .O(N__23471),
            .I(il_min_comp2_D2));
    InMux I__2949 (
            .O(N__23466),
            .I(N__23459));
    InMux I__2948 (
            .O(N__23465),
            .I(N__23459));
    InMux I__2947 (
            .O(N__23464),
            .I(N__23456));
    LocalMux I__2946 (
            .O(N__23459),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__2945 (
            .O(N__23456),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    IoInMux I__2944 (
            .O(N__23451),
            .I(N__23448));
    LocalMux I__2943 (
            .O(N__23448),
            .I(N__23445));
    Span4Mux_s3_v I__2942 (
            .O(N__23445),
            .I(N__23442));
    Span4Mux_v I__2941 (
            .O(N__23442),
            .I(N__23439));
    Span4Mux_v I__2940 (
            .O(N__23439),
            .I(N__23436));
    Span4Mux_v I__2939 (
            .O(N__23436),
            .I(N__23433));
    Odrv4 I__2938 (
            .O(N__23433),
            .I(\delay_measurement_inst.delay_hc_timer.N_393_i ));
    InMux I__2937 (
            .O(N__23430),
            .I(N__23427));
    LocalMux I__2936 (
            .O(N__23427),
            .I(N__23424));
    Span4Mux_h I__2935 (
            .O(N__23424),
            .I(N__23421));
    Odrv4 I__2934 (
            .O(N__23421),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__2933 (
            .O(N__23418),
            .I(N__23415));
    LocalMux I__2932 (
            .O(N__23415),
            .I(N__23411));
    InMux I__2931 (
            .O(N__23414),
            .I(N__23408));
    Odrv4 I__2930 (
            .O(N__23411),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    LocalMux I__2929 (
            .O(N__23408),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    CascadeMux I__2928 (
            .O(N__23403),
            .I(N__23400));
    InMux I__2927 (
            .O(N__23400),
            .I(N__23396));
    InMux I__2926 (
            .O(N__23399),
            .I(N__23393));
    LocalMux I__2925 (
            .O(N__23396),
            .I(N__23388));
    LocalMux I__2924 (
            .O(N__23393),
            .I(N__23388));
    Odrv4 I__2923 (
            .O(N__23388),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2922 (
            .O(N__23385),
            .I(N__23382));
    LocalMux I__2921 (
            .O(N__23382),
            .I(N__23379));
    Span4Mux_h I__2920 (
            .O(N__23379),
            .I(N__23376));
    Odrv4 I__2919 (
            .O(N__23376),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__2918 (
            .O(N__23373),
            .I(N__23370));
    LocalMux I__2917 (
            .O(N__23370),
            .I(N__23367));
    Odrv12 I__2916 (
            .O(N__23367),
            .I(il_min_comp2_D1));
    InMux I__2915 (
            .O(N__23364),
            .I(N__23361));
    LocalMux I__2914 (
            .O(N__23361),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa ));
    InMux I__2913 (
            .O(N__23358),
            .I(N__23355));
    LocalMux I__2912 (
            .O(N__23355),
            .I(N__23352));
    Span4Mux_h I__2911 (
            .O(N__23352),
            .I(N__23349));
    Odrv4 I__2910 (
            .O(N__23349),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__2909 (
            .O(N__23346),
            .I(N__23343));
    LocalMux I__2908 (
            .O(N__23343),
            .I(N__23340));
    Odrv4 I__2907 (
            .O(N__23340),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__2906 (
            .O(N__23337),
            .I(N__23334));
    LocalMux I__2905 (
            .O(N__23334),
            .I(N__23331));
    Odrv4 I__2904 (
            .O(N__23331),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    CascadeMux I__2903 (
            .O(N__23328),
            .I(N__23325));
    InMux I__2902 (
            .O(N__23325),
            .I(N__23322));
    LocalMux I__2901 (
            .O(N__23322),
            .I(N__23319));
    Odrv4 I__2900 (
            .O(N__23319),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__2899 (
            .O(N__23316),
            .I(N__23313));
    LocalMux I__2898 (
            .O(N__23313),
            .I(N__23310));
    Odrv4 I__2897 (
            .O(N__23310),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__2896 (
            .O(N__23307),
            .I(N__23304));
    InMux I__2895 (
            .O(N__23304),
            .I(N__23301));
    LocalMux I__2894 (
            .O(N__23301),
            .I(N__23298));
    Odrv4 I__2893 (
            .O(N__23298),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    InMux I__2892 (
            .O(N__23295),
            .I(N__23292));
    LocalMux I__2891 (
            .O(N__23292),
            .I(N__23289));
    Odrv4 I__2890 (
            .O(N__23289),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__2889 (
            .O(N__23286),
            .I(N__23283));
    LocalMux I__2888 (
            .O(N__23283),
            .I(N__23280));
    Odrv4 I__2887 (
            .O(N__23280),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__2886 (
            .O(N__23277),
            .I(N__23274));
    InMux I__2885 (
            .O(N__23274),
            .I(N__23271));
    LocalMux I__2884 (
            .O(N__23271),
            .I(N__23268));
    Odrv4 I__2883 (
            .O(N__23268),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__2882 (
            .O(N__23265),
            .I(N__23262));
    LocalMux I__2881 (
            .O(N__23262),
            .I(N__23259));
    Span12Mux_v I__2880 (
            .O(N__23259),
            .I(N__23256));
    Odrv12 I__2879 (
            .O(N__23256),
            .I(il_max_comp2_D1));
    InMux I__2878 (
            .O(N__23253),
            .I(N__23250));
    LocalMux I__2877 (
            .O(N__23250),
            .I(N__23247));
    Odrv12 I__2876 (
            .O(N__23247),
            .I(il_min_comp2_c));
    CascadeMux I__2875 (
            .O(N__23244),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__2874 (
            .O(N__23241),
            .I(N__23235));
    InMux I__2873 (
            .O(N__23240),
            .I(N__23235));
    LocalMux I__2872 (
            .O(N__23235),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2871 (
            .O(N__23232),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    CascadeMux I__2870 (
            .O(N__23229),
            .I(N__23225));
    CascadeMux I__2869 (
            .O(N__23228),
            .I(N__23222));
    InMux I__2868 (
            .O(N__23225),
            .I(N__23219));
    InMux I__2867 (
            .O(N__23222),
            .I(N__23216));
    LocalMux I__2866 (
            .O(N__23219),
            .I(N__23211));
    LocalMux I__2865 (
            .O(N__23216),
            .I(N__23211));
    Odrv4 I__2864 (
            .O(N__23211),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2863 (
            .O(N__23208),
            .I(bfn_5_12_0_));
    CascadeMux I__2862 (
            .O(N__23205),
            .I(N__23201));
    InMux I__2861 (
            .O(N__23204),
            .I(N__23198));
    InMux I__2860 (
            .O(N__23201),
            .I(N__23195));
    LocalMux I__2859 (
            .O(N__23198),
            .I(N__23192));
    LocalMux I__2858 (
            .O(N__23195),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    Odrv4 I__2857 (
            .O(N__23192),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2856 (
            .O(N__23187),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    InMux I__2855 (
            .O(N__23184),
            .I(N__23180));
    InMux I__2854 (
            .O(N__23183),
            .I(N__23177));
    LocalMux I__2853 (
            .O(N__23180),
            .I(N__23174));
    LocalMux I__2852 (
            .O(N__23177),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    Odrv4 I__2851 (
            .O(N__23174),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2850 (
            .O(N__23169),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2849 (
            .O(N__23166),
            .I(N__23160));
    InMux I__2848 (
            .O(N__23165),
            .I(N__23160));
    LocalMux I__2847 (
            .O(N__23160),
            .I(N__23157));
    Odrv4 I__2846 (
            .O(N__23157),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2845 (
            .O(N__23154),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2844 (
            .O(N__23151),
            .I(N__23147));
    InMux I__2843 (
            .O(N__23150),
            .I(N__23144));
    LocalMux I__2842 (
            .O(N__23147),
            .I(N__23141));
    LocalMux I__2841 (
            .O(N__23144),
            .I(N__23138));
    Span4Mux_h I__2840 (
            .O(N__23141),
            .I(N__23135));
    Odrv4 I__2839 (
            .O(N__23138),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    Odrv4 I__2838 (
            .O(N__23135),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2837 (
            .O(N__23130),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2836 (
            .O(N__23127),
            .I(N__23121));
    InMux I__2835 (
            .O(N__23126),
            .I(N__23121));
    LocalMux I__2834 (
            .O(N__23121),
            .I(N__23118));
    Odrv4 I__2833 (
            .O(N__23118),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2832 (
            .O(N__23115),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2831 (
            .O(N__23112),
            .I(N__23106));
    InMux I__2830 (
            .O(N__23111),
            .I(N__23106));
    LocalMux I__2829 (
            .O(N__23106),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2828 (
            .O(N__23103),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2827 (
            .O(N__23100),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2826 (
            .O(N__23097),
            .I(N__23091));
    InMux I__2825 (
            .O(N__23096),
            .I(N__23091));
    LocalMux I__2824 (
            .O(N__23091),
            .I(N__23083));
    InMux I__2823 (
            .O(N__23090),
            .I(N__23078));
    InMux I__2822 (
            .O(N__23089),
            .I(N__23078));
    InMux I__2821 (
            .O(N__23088),
            .I(N__23075));
    InMux I__2820 (
            .O(N__23087),
            .I(N__23072));
    InMux I__2819 (
            .O(N__23086),
            .I(N__23069));
    Span4Mux_s2_h I__2818 (
            .O(N__23083),
            .I(N__23055));
    LocalMux I__2817 (
            .O(N__23078),
            .I(N__23055));
    LocalMux I__2816 (
            .O(N__23075),
            .I(N__23055));
    LocalMux I__2815 (
            .O(N__23072),
            .I(N__23055));
    LocalMux I__2814 (
            .O(N__23069),
            .I(N__23055));
    InMux I__2813 (
            .O(N__23068),
            .I(N__23050));
    InMux I__2812 (
            .O(N__23067),
            .I(N__23050));
    InMux I__2811 (
            .O(N__23066),
            .I(N__23047));
    Sp12to4 I__2810 (
            .O(N__23055),
            .I(N__23040));
    LocalMux I__2809 (
            .O(N__23050),
            .I(N__23040));
    LocalMux I__2808 (
            .O(N__23047),
            .I(N__23040));
    Span12Mux_s11_v I__2807 (
            .O(N__23040),
            .I(N__23037));
    Odrv12 I__2806 (
            .O(N__23037),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__2805 (
            .O(N__23034),
            .I(N__23030));
    InMux I__2804 (
            .O(N__23033),
            .I(N__23027));
    LocalMux I__2803 (
            .O(N__23030),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    LocalMux I__2802 (
            .O(N__23027),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2801 (
            .O(N__23022),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    CascadeMux I__2800 (
            .O(N__23019),
            .I(N__23015));
    InMux I__2799 (
            .O(N__23018),
            .I(N__23012));
    InMux I__2798 (
            .O(N__23015),
            .I(N__23009));
    LocalMux I__2797 (
            .O(N__23012),
            .I(N__23006));
    LocalMux I__2796 (
            .O(N__23009),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    Odrv4 I__2795 (
            .O(N__23006),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2794 (
            .O(N__23001),
            .I(bfn_5_11_0_));
    InMux I__2793 (
            .O(N__22998),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    InMux I__2792 (
            .O(N__22995),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    CascadeMux I__2791 (
            .O(N__22992),
            .I(N__22988));
    InMux I__2790 (
            .O(N__22991),
            .I(N__22985));
    InMux I__2789 (
            .O(N__22988),
            .I(N__22982));
    LocalMux I__2788 (
            .O(N__22985),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    LocalMux I__2787 (
            .O(N__22982),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2786 (
            .O(N__22977),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2785 (
            .O(N__22974),
            .I(N__22970));
    InMux I__2784 (
            .O(N__22973),
            .I(N__22967));
    LocalMux I__2783 (
            .O(N__22970),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    LocalMux I__2782 (
            .O(N__22967),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2781 (
            .O(N__22962),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__2780 (
            .O(N__22959),
            .I(N__22955));
    InMux I__2779 (
            .O(N__22958),
            .I(N__22952));
    LocalMux I__2778 (
            .O(N__22955),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__2777 (
            .O(N__22952),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2776 (
            .O(N__22947),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2775 (
            .O(N__22944),
            .I(N__22940));
    InMux I__2774 (
            .O(N__22943),
            .I(N__22937));
    LocalMux I__2773 (
            .O(N__22940),
            .I(N__22934));
    LocalMux I__2772 (
            .O(N__22937),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    Odrv4 I__2771 (
            .O(N__22934),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2770 (
            .O(N__22929),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2769 (
            .O(N__22926),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    CascadeMux I__2768 (
            .O(N__22923),
            .I(N__22920));
    InMux I__2767 (
            .O(N__22920),
            .I(N__22915));
    InMux I__2766 (
            .O(N__22919),
            .I(N__22912));
    InMux I__2765 (
            .O(N__22918),
            .I(N__22909));
    LocalMux I__2764 (
            .O(N__22915),
            .I(N__22906));
    LocalMux I__2763 (
            .O(N__22912),
            .I(N__22901));
    LocalMux I__2762 (
            .O(N__22909),
            .I(N__22901));
    Span4Mux_h I__2761 (
            .O(N__22906),
            .I(N__22898));
    Span12Mux_s8_v I__2760 (
            .O(N__22901),
            .I(N__22895));
    Odrv4 I__2759 (
            .O(N__22898),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv12 I__2758 (
            .O(N__22895),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2757 (
            .O(N__22890),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2756 (
            .O(N__22887),
            .I(N__22882));
    InMux I__2755 (
            .O(N__22886),
            .I(N__22879));
    InMux I__2754 (
            .O(N__22885),
            .I(N__22876));
    LocalMux I__2753 (
            .O(N__22882),
            .I(N__22873));
    LocalMux I__2752 (
            .O(N__22879),
            .I(N__22868));
    LocalMux I__2751 (
            .O(N__22876),
            .I(N__22868));
    Span4Mux_h I__2750 (
            .O(N__22873),
            .I(N__22865));
    Span4Mux_h I__2749 (
            .O(N__22868),
            .I(N__22862));
    Odrv4 I__2748 (
            .O(N__22865),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv4 I__2747 (
            .O(N__22862),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2746 (
            .O(N__22857),
            .I(bfn_5_10_0_));
    InMux I__2745 (
            .O(N__22854),
            .I(N__22850));
    InMux I__2744 (
            .O(N__22853),
            .I(N__22847));
    LocalMux I__2743 (
            .O(N__22850),
            .I(N__22841));
    LocalMux I__2742 (
            .O(N__22847),
            .I(N__22841));
    InMux I__2741 (
            .O(N__22846),
            .I(N__22838));
    Span4Mux_v I__2740 (
            .O(N__22841),
            .I(N__22833));
    LocalMux I__2739 (
            .O(N__22838),
            .I(N__22833));
    Span4Mux_h I__2738 (
            .O(N__22833),
            .I(N__22830));
    Odrv4 I__2737 (
            .O(N__22830),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2736 (
            .O(N__22827),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    InMux I__2735 (
            .O(N__22824),
            .I(N__22818));
    InMux I__2734 (
            .O(N__22823),
            .I(N__22818));
    LocalMux I__2733 (
            .O(N__22818),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2732 (
            .O(N__22815),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2731 (
            .O(N__22812),
            .I(N__22806));
    InMux I__2730 (
            .O(N__22811),
            .I(N__22806));
    LocalMux I__2729 (
            .O(N__22806),
            .I(N__22803));
    Odrv4 I__2728 (
            .O(N__22803),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2727 (
            .O(N__22800),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    CascadeMux I__2726 (
            .O(N__22797),
            .I(N__22794));
    InMux I__2725 (
            .O(N__22794),
            .I(N__22788));
    InMux I__2724 (
            .O(N__22793),
            .I(N__22788));
    LocalMux I__2723 (
            .O(N__22788),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2722 (
            .O(N__22785),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2721 (
            .O(N__22782),
            .I(N__22776));
    InMux I__2720 (
            .O(N__22781),
            .I(N__22776));
    LocalMux I__2719 (
            .O(N__22776),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2718 (
            .O(N__22773),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2717 (
            .O(N__22770),
            .I(N__22764));
    InMux I__2716 (
            .O(N__22769),
            .I(N__22764));
    LocalMux I__2715 (
            .O(N__22764),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2714 (
            .O(N__22761),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2713 (
            .O(N__22758),
            .I(N__22755));
    LocalMux I__2712 (
            .O(N__22755),
            .I(N__22752));
    Span4Mux_h I__2711 (
            .O(N__22752),
            .I(N__22749));
    Odrv4 I__2710 (
            .O(N__22749),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2709 (
            .O(N__22746),
            .I(N__22743));
    LocalMux I__2708 (
            .O(N__22743),
            .I(N__22740));
    Odrv12 I__2707 (
            .O(N__22740),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__2706 (
            .O(N__22737),
            .I(N__22734));
    LocalMux I__2705 (
            .O(N__22734),
            .I(N__22731));
    Span4Mux_h I__2704 (
            .O(N__22731),
            .I(N__22728));
    Odrv4 I__2703 (
            .O(N__22728),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2702 (
            .O(N__22725),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    InMux I__2701 (
            .O(N__22722),
            .I(N__22719));
    LocalMux I__2700 (
            .O(N__22719),
            .I(N__22716));
    Span4Mux_h I__2699 (
            .O(N__22716),
            .I(N__22713));
    Odrv4 I__2698 (
            .O(N__22713),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2697 (
            .O(N__22710),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2696 (
            .O(N__22707),
            .I(N__22704));
    LocalMux I__2695 (
            .O(N__22704),
            .I(N__22699));
    InMux I__2694 (
            .O(N__22703),
            .I(N__22696));
    InMux I__2693 (
            .O(N__22702),
            .I(N__22693));
    Span4Mux_s2_h I__2692 (
            .O(N__22699),
            .I(N__22688));
    LocalMux I__2691 (
            .O(N__22696),
            .I(N__22688));
    LocalMux I__2690 (
            .O(N__22693),
            .I(N__22685));
    Span4Mux_h I__2689 (
            .O(N__22688),
            .I(N__22682));
    Span4Mux_h I__2688 (
            .O(N__22685),
            .I(N__22679));
    Odrv4 I__2687 (
            .O(N__22682),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__2686 (
            .O(N__22679),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2685 (
            .O(N__22674),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    CascadeMux I__2684 (
            .O(N__22671),
            .I(N__22668));
    InMux I__2683 (
            .O(N__22668),
            .I(N__22665));
    LocalMux I__2682 (
            .O(N__22665),
            .I(N__22661));
    InMux I__2681 (
            .O(N__22664),
            .I(N__22658));
    Span4Mux_v I__2680 (
            .O(N__22661),
            .I(N__22651));
    LocalMux I__2679 (
            .O(N__22658),
            .I(N__22651));
    InMux I__2678 (
            .O(N__22657),
            .I(N__22646));
    InMux I__2677 (
            .O(N__22656),
            .I(N__22646));
    Span4Mux_s2_h I__2676 (
            .O(N__22651),
            .I(N__22641));
    LocalMux I__2675 (
            .O(N__22646),
            .I(N__22641));
    Span4Mux_h I__2674 (
            .O(N__22641),
            .I(N__22638));
    Odrv4 I__2673 (
            .O(N__22638),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2672 (
            .O(N__22635),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    CascadeMux I__2671 (
            .O(N__22632),
            .I(N__22629));
    InMux I__2670 (
            .O(N__22629),
            .I(N__22626));
    LocalMux I__2669 (
            .O(N__22626),
            .I(N__22621));
    InMux I__2668 (
            .O(N__22625),
            .I(N__22618));
    InMux I__2667 (
            .O(N__22624),
            .I(N__22615));
    Span4Mux_v I__2666 (
            .O(N__22621),
            .I(N__22610));
    LocalMux I__2665 (
            .O(N__22618),
            .I(N__22610));
    LocalMux I__2664 (
            .O(N__22615),
            .I(N__22607));
    Span4Mux_h I__2663 (
            .O(N__22610),
            .I(N__22604));
    Span4Mux_h I__2662 (
            .O(N__22607),
            .I(N__22601));
    Odrv4 I__2661 (
            .O(N__22604),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__2660 (
            .O(N__22601),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2659 (
            .O(N__22596),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    CascadeMux I__2658 (
            .O(N__22593),
            .I(N__22590));
    InMux I__2657 (
            .O(N__22590),
            .I(N__22586));
    InMux I__2656 (
            .O(N__22589),
            .I(N__22582));
    LocalMux I__2655 (
            .O(N__22586),
            .I(N__22579));
    InMux I__2654 (
            .O(N__22585),
            .I(N__22576));
    LocalMux I__2653 (
            .O(N__22582),
            .I(N__22573));
    Span4Mux_v I__2652 (
            .O(N__22579),
            .I(N__22568));
    LocalMux I__2651 (
            .O(N__22576),
            .I(N__22568));
    Span4Mux_h I__2650 (
            .O(N__22573),
            .I(N__22565));
    Span4Mux_h I__2649 (
            .O(N__22568),
            .I(N__22562));
    Odrv4 I__2648 (
            .O(N__22565),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2647 (
            .O(N__22562),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2646 (
            .O(N__22557),
            .I(N__22552));
    InMux I__2645 (
            .O(N__22556),
            .I(N__22549));
    InMux I__2644 (
            .O(N__22555),
            .I(N__22546));
    LocalMux I__2643 (
            .O(N__22552),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2642 (
            .O(N__22549),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2641 (
            .O(N__22546),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__2640 (
            .O(N__22539),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__2639 (
            .O(N__22536),
            .I(N__22531));
    InMux I__2638 (
            .O(N__22535),
            .I(N__22528));
    InMux I__2637 (
            .O(N__22534),
            .I(N__22525));
    LocalMux I__2636 (
            .O(N__22531),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2635 (
            .O(N__22528),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2634 (
            .O(N__22525),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2633 (
            .O(N__22518),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__2632 (
            .O(N__22515),
            .I(N__22510));
    InMux I__2631 (
            .O(N__22514),
            .I(N__22507));
    InMux I__2630 (
            .O(N__22513),
            .I(N__22504));
    LocalMux I__2629 (
            .O(N__22510),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2628 (
            .O(N__22507),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2627 (
            .O(N__22504),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__2626 (
            .O(N__22497),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__2625 (
            .O(N__22494),
            .I(N__22489));
    InMux I__2624 (
            .O(N__22493),
            .I(N__22486));
    InMux I__2623 (
            .O(N__22492),
            .I(N__22483));
    LocalMux I__2622 (
            .O(N__22489),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2621 (
            .O(N__22486),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2620 (
            .O(N__22483),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__2619 (
            .O(N__22476),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__2618 (
            .O(N__22473),
            .I(N__22468));
    InMux I__2617 (
            .O(N__22472),
            .I(N__22465));
    InMux I__2616 (
            .O(N__22471),
            .I(N__22462));
    LocalMux I__2615 (
            .O(N__22468),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2614 (
            .O(N__22465),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2613 (
            .O(N__22462),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2612 (
            .O(N__22455),
            .I(bfn_4_13_0_));
    InMux I__2611 (
            .O(N__22452),
            .I(N__22434));
    InMux I__2610 (
            .O(N__22451),
            .I(N__22434));
    InMux I__2609 (
            .O(N__22450),
            .I(N__22434));
    InMux I__2608 (
            .O(N__22449),
            .I(N__22434));
    InMux I__2607 (
            .O(N__22448),
            .I(N__22429));
    InMux I__2606 (
            .O(N__22447),
            .I(N__22429));
    InMux I__2605 (
            .O(N__22446),
            .I(N__22420));
    InMux I__2604 (
            .O(N__22445),
            .I(N__22420));
    InMux I__2603 (
            .O(N__22444),
            .I(N__22420));
    InMux I__2602 (
            .O(N__22443),
            .I(N__22420));
    LocalMux I__2601 (
            .O(N__22434),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__2600 (
            .O(N__22429),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__2599 (
            .O(N__22420),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__2598 (
            .O(N__22413),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__2597 (
            .O(N__22410),
            .I(N__22405));
    InMux I__2596 (
            .O(N__22409),
            .I(N__22402));
    InMux I__2595 (
            .O(N__22408),
            .I(N__22399));
    LocalMux I__2594 (
            .O(N__22405),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2593 (
            .O(N__22402),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2592 (
            .O(N__22399),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    CascadeMux I__2591 (
            .O(N__22392),
            .I(N__22389));
    InMux I__2590 (
            .O(N__22389),
            .I(N__22386));
    LocalMux I__2589 (
            .O(N__22386),
            .I(N__22382));
    InMux I__2588 (
            .O(N__22385),
            .I(N__22379));
    Span4Mux_h I__2587 (
            .O(N__22382),
            .I(N__22374));
    LocalMux I__2586 (
            .O(N__22379),
            .I(N__22374));
    Span4Mux_v I__2585 (
            .O(N__22374),
            .I(N__22371));
    Span4Mux_h I__2584 (
            .O(N__22371),
            .I(N__22368));
    Span4Mux_v I__2583 (
            .O(N__22368),
            .I(N__22365));
    Odrv4 I__2582 (
            .O(N__22365),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__2581 (
            .O(N__22362),
            .I(N__22358));
    InMux I__2580 (
            .O(N__22361),
            .I(N__22354));
    LocalMux I__2579 (
            .O(N__22358),
            .I(N__22351));
    InMux I__2578 (
            .O(N__22357),
            .I(N__22348));
    LocalMux I__2577 (
            .O(N__22354),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    Odrv12 I__2576 (
            .O(N__22351),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    LocalMux I__2575 (
            .O(N__22348),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ));
    InMux I__2574 (
            .O(N__22341),
            .I(N__22338));
    LocalMux I__2573 (
            .O(N__22338),
            .I(N__22335));
    Odrv12 I__2572 (
            .O(N__22335),
            .I(il_max_comp2_c));
    InMux I__2571 (
            .O(N__22332),
            .I(N__22329));
    LocalMux I__2570 (
            .O(N__22329),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__2569 (
            .O(N__22326),
            .I(N__22323));
    InMux I__2568 (
            .O(N__22323),
            .I(N__22320));
    LocalMux I__2567 (
            .O(N__22320),
            .I(N__22317));
    Odrv4 I__2566 (
            .O(N__22317),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__2565 (
            .O(N__22314),
            .I(N__22311));
    LocalMux I__2564 (
            .O(N__22311),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    CascadeMux I__2563 (
            .O(N__22308),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ));
    InMux I__2562 (
            .O(N__22305),
            .I(N__22302));
    LocalMux I__2561 (
            .O(N__22302),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2560 (
            .O(N__22299),
            .I(N__22294));
    InMux I__2559 (
            .O(N__22298),
            .I(N__22291));
    InMux I__2558 (
            .O(N__22297),
            .I(N__22288));
    LocalMux I__2557 (
            .O(N__22294),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2556 (
            .O(N__22291),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2555 (
            .O(N__22288),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2554 (
            .O(N__22281),
            .I(bfn_4_12_0_));
    InMux I__2553 (
            .O(N__22278),
            .I(N__22273));
    InMux I__2552 (
            .O(N__22277),
            .I(N__22270));
    InMux I__2551 (
            .O(N__22276),
            .I(N__22267));
    LocalMux I__2550 (
            .O(N__22273),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2549 (
            .O(N__22270),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2548 (
            .O(N__22267),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__2547 (
            .O(N__22260),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__2546 (
            .O(N__22257),
            .I(N__22252));
    InMux I__2545 (
            .O(N__22256),
            .I(N__22249));
    InMux I__2544 (
            .O(N__22255),
            .I(N__22246));
    LocalMux I__2543 (
            .O(N__22252),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2542 (
            .O(N__22249),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2541 (
            .O(N__22246),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2540 (
            .O(N__22239),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__2539 (
            .O(N__22236),
            .I(N__22231));
    InMux I__2538 (
            .O(N__22235),
            .I(N__22228));
    InMux I__2537 (
            .O(N__22234),
            .I(N__22225));
    LocalMux I__2536 (
            .O(N__22231),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2535 (
            .O(N__22228),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2534 (
            .O(N__22225),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__2533 (
            .O(N__22218),
            .I(\pwm_generator_inst.counter_cry_2 ));
    CascadeMux I__2532 (
            .O(N__22215),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    InMux I__2531 (
            .O(N__22212),
            .I(N__22209));
    LocalMux I__2530 (
            .O(N__22209),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    CascadeMux I__2529 (
            .O(N__22206),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ));
    InMux I__2528 (
            .O(N__22203),
            .I(N__22195));
    InMux I__2527 (
            .O(N__22202),
            .I(N__22195));
    CascadeMux I__2526 (
            .O(N__22201),
            .I(N__22190));
    CascadeMux I__2525 (
            .O(N__22200),
            .I(N__22187));
    LocalMux I__2524 (
            .O(N__22195),
            .I(N__22181));
    InMux I__2523 (
            .O(N__22194),
            .I(N__22174));
    InMux I__2522 (
            .O(N__22193),
            .I(N__22174));
    InMux I__2521 (
            .O(N__22190),
            .I(N__22174));
    InMux I__2520 (
            .O(N__22187),
            .I(N__22171));
    InMux I__2519 (
            .O(N__22186),
            .I(N__22168));
    InMux I__2518 (
            .O(N__22185),
            .I(N__22165));
    InMux I__2517 (
            .O(N__22184),
            .I(N__22162));
    Span4Mux_v I__2516 (
            .O(N__22181),
            .I(N__22159));
    LocalMux I__2515 (
            .O(N__22174),
            .I(N__22154));
    LocalMux I__2514 (
            .O(N__22171),
            .I(N__22154));
    LocalMux I__2513 (
            .O(N__22168),
            .I(N__22151));
    LocalMux I__2512 (
            .O(N__22165),
            .I(N__22146));
    LocalMux I__2511 (
            .O(N__22162),
            .I(N__22146));
    Span4Mux_h I__2510 (
            .O(N__22159),
            .I(N__22143));
    Span4Mux_h I__2509 (
            .O(N__22154),
            .I(N__22140));
    Span4Mux_h I__2508 (
            .O(N__22151),
            .I(N__22137));
    Span4Mux_h I__2507 (
            .O(N__22146),
            .I(N__22134));
    Odrv4 I__2506 (
            .O(N__22143),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2505 (
            .O(N__22140),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2504 (
            .O(N__22137),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2503 (
            .O(N__22134),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    InMux I__2502 (
            .O(N__22125),
            .I(N__22122));
    LocalMux I__2501 (
            .O(N__22122),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    CascadeMux I__2500 (
            .O(N__22119),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ));
    InMux I__2499 (
            .O(N__22116),
            .I(N__22113));
    LocalMux I__2498 (
            .O(N__22113),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    InMux I__2497 (
            .O(N__22110),
            .I(N__22107));
    LocalMux I__2496 (
            .O(N__22107),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__2495 (
            .O(N__22104),
            .I(N__22101));
    LocalMux I__2494 (
            .O(N__22101),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__2493 (
            .O(N__22098),
            .I(N__22095));
    LocalMux I__2492 (
            .O(N__22095),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ));
    InMux I__2491 (
            .O(N__22092),
            .I(N__22089));
    LocalMux I__2490 (
            .O(N__22089),
            .I(N__22086));
    Odrv12 I__2489 (
            .O(N__22086),
            .I(\pwm_generator_inst.thresholdZ0Z_5 ));
    InMux I__2488 (
            .O(N__22083),
            .I(N__22080));
    LocalMux I__2487 (
            .O(N__22080),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_0 ));
    InMux I__2486 (
            .O(N__22077),
            .I(N__22074));
    LocalMux I__2485 (
            .O(N__22074),
            .I(N__22071));
    Span12Mux_s11_v I__2484 (
            .O(N__22071),
            .I(N__22068));
    Odrv12 I__2483 (
            .O(N__22068),
            .I(\pwm_generator_inst.thresholdZ0Z_0 ));
    InMux I__2482 (
            .O(N__22065),
            .I(N__22062));
    LocalMux I__2481 (
            .O(N__22062),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ));
    InMux I__2480 (
            .O(N__22059),
            .I(N__22056));
    LocalMux I__2479 (
            .O(N__22056),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_5 ));
    CascadeMux I__2478 (
            .O(N__22053),
            .I(N__22050));
    InMux I__2477 (
            .O(N__22050),
            .I(N__22047));
    LocalMux I__2476 (
            .O(N__22047),
            .I(N__22044));
    Odrv12 I__2475 (
            .O(N__22044),
            .I(\pwm_generator_inst.thresholdZ0Z_9 ));
    InMux I__2474 (
            .O(N__22041),
            .I(N__22038));
    LocalMux I__2473 (
            .O(N__22038),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ));
    InMux I__2472 (
            .O(N__22035),
            .I(N__22032));
    LocalMux I__2471 (
            .O(N__22032),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_9 ));
    InMux I__2470 (
            .O(N__22029),
            .I(N__22026));
    LocalMux I__2469 (
            .O(N__22026),
            .I(N__22023));
    Odrv12 I__2468 (
            .O(N__22023),
            .I(\pwm_generator_inst.thresholdZ0Z_8 ));
    InMux I__2467 (
            .O(N__22020),
            .I(N__22013));
    InMux I__2466 (
            .O(N__22019),
            .I(N__22013));
    InMux I__2465 (
            .O(N__22018),
            .I(N__22010));
    LocalMux I__2464 (
            .O(N__22013),
            .I(N__22005));
    LocalMux I__2463 (
            .O(N__22010),
            .I(N__22002));
    InMux I__2462 (
            .O(N__22009),
            .I(N__21997));
    InMux I__2461 (
            .O(N__22008),
            .I(N__21997));
    Span4Mux_v I__2460 (
            .O(N__22005),
            .I(N__21990));
    Span4Mux_s3_h I__2459 (
            .O(N__22002),
            .I(N__21990));
    LocalMux I__2458 (
            .O(N__21997),
            .I(N__21990));
    Span4Mux_v I__2457 (
            .O(N__21990),
            .I(N__21982));
    InMux I__2456 (
            .O(N__21989),
            .I(N__21979));
    InMux I__2455 (
            .O(N__21988),
            .I(N__21976));
    InMux I__2454 (
            .O(N__21987),
            .I(N__21969));
    InMux I__2453 (
            .O(N__21986),
            .I(N__21969));
    InMux I__2452 (
            .O(N__21985),
            .I(N__21969));
    Span4Mux_v I__2451 (
            .O(N__21982),
            .I(N__21966));
    LocalMux I__2450 (
            .O(N__21979),
            .I(N__21961));
    LocalMux I__2449 (
            .O(N__21976),
            .I(N__21961));
    LocalMux I__2448 (
            .O(N__21969),
            .I(N__21958));
    Odrv4 I__2447 (
            .O(N__21966),
            .I(\pwm_generator_inst.N_16 ));
    Odrv12 I__2446 (
            .O(N__21961),
            .I(\pwm_generator_inst.N_16 ));
    Odrv4 I__2445 (
            .O(N__21958),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__2444 (
            .O(N__21951),
            .I(N__21944));
    CascadeMux I__2443 (
            .O(N__21950),
            .I(N__21940));
    CascadeMux I__2442 (
            .O(N__21949),
            .I(N__21936));
    CascadeMux I__2441 (
            .O(N__21948),
            .I(N__21933));
    InMux I__2440 (
            .O(N__21947),
            .I(N__21928));
    InMux I__2439 (
            .O(N__21944),
            .I(N__21928));
    InMux I__2438 (
            .O(N__21943),
            .I(N__21908));
    InMux I__2437 (
            .O(N__21940),
            .I(N__21905));
    CascadeMux I__2436 (
            .O(N__21939),
            .I(N__21902));
    InMux I__2435 (
            .O(N__21936),
            .I(N__21897));
    InMux I__2434 (
            .O(N__21933),
            .I(N__21897));
    LocalMux I__2433 (
            .O(N__21928),
            .I(N__21894));
    InMux I__2432 (
            .O(N__21927),
            .I(N__21888));
    InMux I__2431 (
            .O(N__21926),
            .I(N__21871));
    InMux I__2430 (
            .O(N__21925),
            .I(N__21871));
    InMux I__2429 (
            .O(N__21924),
            .I(N__21871));
    InMux I__2428 (
            .O(N__21923),
            .I(N__21871));
    InMux I__2427 (
            .O(N__21922),
            .I(N__21871));
    InMux I__2426 (
            .O(N__21921),
            .I(N__21871));
    InMux I__2425 (
            .O(N__21920),
            .I(N__21871));
    InMux I__2424 (
            .O(N__21919),
            .I(N__21871));
    InMux I__2423 (
            .O(N__21918),
            .I(N__21856));
    InMux I__2422 (
            .O(N__21917),
            .I(N__21856));
    InMux I__2421 (
            .O(N__21916),
            .I(N__21856));
    InMux I__2420 (
            .O(N__21915),
            .I(N__21856));
    InMux I__2419 (
            .O(N__21914),
            .I(N__21856));
    InMux I__2418 (
            .O(N__21913),
            .I(N__21856));
    InMux I__2417 (
            .O(N__21912),
            .I(N__21856));
    CascadeMux I__2416 (
            .O(N__21911),
            .I(N__21848));
    LocalMux I__2415 (
            .O(N__21908),
            .I(N__21843));
    LocalMux I__2414 (
            .O(N__21905),
            .I(N__21843));
    InMux I__2413 (
            .O(N__21902),
            .I(N__21840));
    LocalMux I__2412 (
            .O(N__21897),
            .I(N__21837));
    Span4Mux_h I__2411 (
            .O(N__21894),
            .I(N__21834));
    CascadeMux I__2410 (
            .O(N__21893),
            .I(N__21831));
    InMux I__2409 (
            .O(N__21892),
            .I(N__21826));
    InMux I__2408 (
            .O(N__21891),
            .I(N__21826));
    LocalMux I__2407 (
            .O(N__21888),
            .I(N__21819));
    LocalMux I__2406 (
            .O(N__21871),
            .I(N__21819));
    LocalMux I__2405 (
            .O(N__21856),
            .I(N__21819));
    InMux I__2404 (
            .O(N__21855),
            .I(N__21812));
    InMux I__2403 (
            .O(N__21854),
            .I(N__21812));
    InMux I__2402 (
            .O(N__21853),
            .I(N__21812));
    InMux I__2401 (
            .O(N__21852),
            .I(N__21805));
    InMux I__2400 (
            .O(N__21851),
            .I(N__21805));
    InMux I__2399 (
            .O(N__21848),
            .I(N__21805));
    Span4Mux_v I__2398 (
            .O(N__21843),
            .I(N__21802));
    LocalMux I__2397 (
            .O(N__21840),
            .I(N__21795));
    Span12Mux_h I__2396 (
            .O(N__21837),
            .I(N__21795));
    Sp12to4 I__2395 (
            .O(N__21834),
            .I(N__21795));
    InMux I__2394 (
            .O(N__21831),
            .I(N__21792));
    LocalMux I__2393 (
            .O(N__21826),
            .I(N__21789));
    Span4Mux_v I__2392 (
            .O(N__21819),
            .I(N__21784));
    LocalMux I__2391 (
            .O(N__21812),
            .I(N__21784));
    LocalMux I__2390 (
            .O(N__21805),
            .I(N_19_1));
    Odrv4 I__2389 (
            .O(N__21802),
            .I(N_19_1));
    Odrv12 I__2388 (
            .O(N__21795),
            .I(N_19_1));
    LocalMux I__2387 (
            .O(N__21792),
            .I(N_19_1));
    Odrv4 I__2386 (
            .O(N__21789),
            .I(N_19_1));
    Odrv4 I__2385 (
            .O(N__21784),
            .I(N_19_1));
    CascadeMux I__2384 (
            .O(N__21771),
            .I(N__21768));
    InMux I__2383 (
            .O(N__21768),
            .I(N__21765));
    LocalMux I__2382 (
            .O(N__21765),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ));
    InMux I__2381 (
            .O(N__21762),
            .I(N__21753));
    InMux I__2380 (
            .O(N__21761),
            .I(N__21753));
    InMux I__2379 (
            .O(N__21760),
            .I(N__21748));
    InMux I__2378 (
            .O(N__21759),
            .I(N__21748));
    InMux I__2377 (
            .O(N__21758),
            .I(N__21745));
    LocalMux I__2376 (
            .O(N__21753),
            .I(N__21742));
    LocalMux I__2375 (
            .O(N__21748),
            .I(N__21737));
    LocalMux I__2374 (
            .O(N__21745),
            .I(N__21732));
    Span4Mux_h I__2373 (
            .O(N__21742),
            .I(N__21732));
    InMux I__2372 (
            .O(N__21741),
            .I(N__21729));
    InMux I__2371 (
            .O(N__21740),
            .I(N__21726));
    Span12Mux_s6_h I__2370 (
            .O(N__21737),
            .I(N__21720));
    Span4Mux_v I__2369 (
            .O(N__21732),
            .I(N__21713));
    LocalMux I__2368 (
            .O(N__21729),
            .I(N__21713));
    LocalMux I__2367 (
            .O(N__21726),
            .I(N__21713));
    InMux I__2366 (
            .O(N__21725),
            .I(N__21706));
    InMux I__2365 (
            .O(N__21724),
            .I(N__21706));
    InMux I__2364 (
            .O(N__21723),
            .I(N__21706));
    Span12Mux_v I__2363 (
            .O(N__21720),
            .I(N__21703));
    Span4Mux_v I__2362 (
            .O(N__21713),
            .I(N__21698));
    LocalMux I__2361 (
            .O(N__21706),
            .I(N__21698));
    Odrv12 I__2360 (
            .O(N__21703),
            .I(\pwm_generator_inst.N_17 ));
    Odrv4 I__2359 (
            .O(N__21698),
            .I(\pwm_generator_inst.N_17 ));
    InMux I__2358 (
            .O(N__21693),
            .I(N__21690));
    LocalMux I__2357 (
            .O(N__21690),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_8 ));
    InMux I__2356 (
            .O(N__21687),
            .I(N__21682));
    InMux I__2355 (
            .O(N__21686),
            .I(N__21679));
    InMux I__2354 (
            .O(N__21685),
            .I(N__21676));
    LocalMux I__2353 (
            .O(N__21682),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__2352 (
            .O(N__21679),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    LocalMux I__2351 (
            .O(N__21676),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ));
    InMux I__2350 (
            .O(N__21669),
            .I(N__21666));
    LocalMux I__2349 (
            .O(N__21666),
            .I(N__21663));
    Span4Mux_v I__2348 (
            .O(N__21663),
            .I(N__21660));
    Odrv4 I__2347 (
            .O(N__21660),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ));
    InMux I__2346 (
            .O(N__21657),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ));
    InMux I__2345 (
            .O(N__21654),
            .I(N__21650));
    InMux I__2344 (
            .O(N__21653),
            .I(N__21646));
    LocalMux I__2343 (
            .O(N__21650),
            .I(N__21643));
    InMux I__2342 (
            .O(N__21649),
            .I(N__21640));
    LocalMux I__2341 (
            .O(N__21646),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    Odrv4 I__2340 (
            .O(N__21643),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    LocalMux I__2339 (
            .O(N__21640),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ));
    InMux I__2338 (
            .O(N__21633),
            .I(N__21630));
    LocalMux I__2337 (
            .O(N__21630),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ));
    InMux I__2336 (
            .O(N__21627),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ));
    InMux I__2335 (
            .O(N__21624),
            .I(N__21621));
    LocalMux I__2334 (
            .O(N__21621),
            .I(N__21616));
    InMux I__2333 (
            .O(N__21620),
            .I(N__21613));
    InMux I__2332 (
            .O(N__21619),
            .I(N__21610));
    Span4Mux_s3_h I__2331 (
            .O(N__21616),
            .I(N__21605));
    LocalMux I__2330 (
            .O(N__21613),
            .I(N__21605));
    LocalMux I__2329 (
            .O(N__21610),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    Odrv4 I__2328 (
            .O(N__21605),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ));
    InMux I__2327 (
            .O(N__21600),
            .I(N__21597));
    LocalMux I__2326 (
            .O(N__21597),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ));
    InMux I__2325 (
            .O(N__21594),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ));
    InMux I__2324 (
            .O(N__21591),
            .I(N__21587));
    InMux I__2323 (
            .O(N__21590),
            .I(N__21584));
    LocalMux I__2322 (
            .O(N__21587),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    LocalMux I__2321 (
            .O(N__21584),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ));
    InMux I__2320 (
            .O(N__21579),
            .I(N__21576));
    LocalMux I__2319 (
            .O(N__21576),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ));
    InMux I__2318 (
            .O(N__21573),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ));
    InMux I__2317 (
            .O(N__21570),
            .I(N__21566));
    InMux I__2316 (
            .O(N__21569),
            .I(N__21563));
    LocalMux I__2315 (
            .O(N__21566),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    LocalMux I__2314 (
            .O(N__21563),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ));
    InMux I__2313 (
            .O(N__21558),
            .I(N__21555));
    LocalMux I__2312 (
            .O(N__21555),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ));
    InMux I__2311 (
            .O(N__21552),
            .I(bfn_3_17_0_));
    InMux I__2310 (
            .O(N__21549),
            .I(N__21545));
    InMux I__2309 (
            .O(N__21548),
            .I(N__21542));
    LocalMux I__2308 (
            .O(N__21545),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    LocalMux I__2307 (
            .O(N__21542),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ));
    InMux I__2306 (
            .O(N__21537),
            .I(N__21534));
    LocalMux I__2305 (
            .O(N__21534),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ));
    InMux I__2304 (
            .O(N__21531),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ));
    InMux I__2303 (
            .O(N__21528),
            .I(N__21523));
    InMux I__2302 (
            .O(N__21527),
            .I(N__21520));
    InMux I__2301 (
            .O(N__21526),
            .I(N__21517));
    LocalMux I__2300 (
            .O(N__21523),
            .I(N__21514));
    LocalMux I__2299 (
            .O(N__21520),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    LocalMux I__2298 (
            .O(N__21517),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    Odrv4 I__2297 (
            .O(N__21514),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ));
    InMux I__2296 (
            .O(N__21507),
            .I(N__21504));
    LocalMux I__2295 (
            .O(N__21504),
            .I(N__21501));
    Odrv4 I__2294 (
            .O(N__21501),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ));
    InMux I__2293 (
            .O(N__21498),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ));
    InMux I__2292 (
            .O(N__21495),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ));
    InMux I__2291 (
            .O(N__21492),
            .I(N__21489));
    LocalMux I__2290 (
            .O(N__21489),
            .I(N__21486));
    Odrv4 I__2289 (
            .O(N__21486),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ));
    InMux I__2288 (
            .O(N__21483),
            .I(N__21480));
    LocalMux I__2287 (
            .O(N__21480),
            .I(N__21477));
    Sp12to4 I__2286 (
            .O(N__21477),
            .I(N__21474));
    Span12Mux_v I__2285 (
            .O(N__21474),
            .I(N__21471));
    Odrv12 I__2284 (
            .O(N__21471),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__2283 (
            .O(N__21468),
            .I(N__21465));
    LocalMux I__2282 (
            .O(N__21465),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ));
    InMux I__2281 (
            .O(N__21462),
            .I(N__21459));
    LocalMux I__2280 (
            .O(N__21459),
            .I(N__21456));
    Span12Mux_v I__2279 (
            .O(N__21456),
            .I(N__21453));
    Odrv12 I__2278 (
            .O(N__21453),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__2277 (
            .O(N__21450),
            .I(N__21447));
    LocalMux I__2276 (
            .O(N__21447),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ));
    InMux I__2275 (
            .O(N__21444),
            .I(N__21441));
    LocalMux I__2274 (
            .O(N__21441),
            .I(N__21438));
    Span4Mux_v I__2273 (
            .O(N__21438),
            .I(N__21435));
    Span4Mux_h I__2272 (
            .O(N__21435),
            .I(N__21432));
    Span4Mux_v I__2271 (
            .O(N__21432),
            .I(N__21429));
    Odrv4 I__2270 (
            .O(N__21429),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__2269 (
            .O(N__21426),
            .I(N__21423));
    LocalMux I__2268 (
            .O(N__21423),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ));
    InMux I__2267 (
            .O(N__21420),
            .I(N__21417));
    LocalMux I__2266 (
            .O(N__21417),
            .I(N__21414));
    Span4Mux_v I__2265 (
            .O(N__21414),
            .I(N__21411));
    Span4Mux_h I__2264 (
            .O(N__21411),
            .I(N__21408));
    Span4Mux_v I__2263 (
            .O(N__21408),
            .I(N__21405));
    Odrv4 I__2262 (
            .O(N__21405),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__2261 (
            .O(N__21402),
            .I(N__21399));
    LocalMux I__2260 (
            .O(N__21399),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ));
    InMux I__2259 (
            .O(N__21396),
            .I(N__21393));
    LocalMux I__2258 (
            .O(N__21393),
            .I(N__21390));
    Span4Mux_h I__2257 (
            .O(N__21390),
            .I(N__21387));
    Span4Mux_v I__2256 (
            .O(N__21387),
            .I(N__21384));
    Span4Mux_v I__2255 (
            .O(N__21384),
            .I(N__21381));
    Odrv4 I__2254 (
            .O(N__21381),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__2253 (
            .O(N__21378),
            .I(N__21375));
    LocalMux I__2252 (
            .O(N__21375),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ));
    InMux I__2251 (
            .O(N__21372),
            .I(N__21369));
    LocalMux I__2250 (
            .O(N__21369),
            .I(N__21366));
    Span4Mux_h I__2249 (
            .O(N__21366),
            .I(N__21363));
    Sp12to4 I__2248 (
            .O(N__21363),
            .I(N__21360));
    Odrv12 I__2247 (
            .O(N__21360),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__2246 (
            .O(N__21357),
            .I(N__21354));
    LocalMux I__2245 (
            .O(N__21354),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ));
    InMux I__2244 (
            .O(N__21351),
            .I(N__21348));
    LocalMux I__2243 (
            .O(N__21348),
            .I(N__21345));
    Span4Mux_s3_h I__2242 (
            .O(N__21345),
            .I(N__21342));
    Odrv4 I__2241 (
            .O(N__21342),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ));
    InMux I__2240 (
            .O(N__21339),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ));
    CascadeMux I__2239 (
            .O(N__21336),
            .I(N__21332));
    CascadeMux I__2238 (
            .O(N__21335),
            .I(N__21328));
    InMux I__2237 (
            .O(N__21332),
            .I(N__21324));
    InMux I__2236 (
            .O(N__21331),
            .I(N__21319));
    InMux I__2235 (
            .O(N__21328),
            .I(N__21316));
    InMux I__2234 (
            .O(N__21327),
            .I(N__21313));
    LocalMux I__2233 (
            .O(N__21324),
            .I(N__21309));
    InMux I__2232 (
            .O(N__21323),
            .I(N__21304));
    InMux I__2231 (
            .O(N__21322),
            .I(N__21304));
    LocalMux I__2230 (
            .O(N__21319),
            .I(N__21297));
    LocalMux I__2229 (
            .O(N__21316),
            .I(N__21297));
    LocalMux I__2228 (
            .O(N__21313),
            .I(N__21297));
    InMux I__2227 (
            .O(N__21312),
            .I(N__21289));
    Span4Mux_v I__2226 (
            .O(N__21309),
            .I(N__21284));
    LocalMux I__2225 (
            .O(N__21304),
            .I(N__21284));
    Span4Mux_v I__2224 (
            .O(N__21297),
            .I(N__21281));
    InMux I__2223 (
            .O(N__21296),
            .I(N__21274));
    InMux I__2222 (
            .O(N__21295),
            .I(N__21274));
    InMux I__2221 (
            .O(N__21294),
            .I(N__21274));
    InMux I__2220 (
            .O(N__21293),
            .I(N__21269));
    InMux I__2219 (
            .O(N__21292),
            .I(N__21269));
    LocalMux I__2218 (
            .O(N__21289),
            .I(N__21266));
    Odrv4 I__2217 (
            .O(N__21284),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv4 I__2216 (
            .O(N__21281),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2215 (
            .O(N__21274),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    LocalMux I__2214 (
            .O(N__21269),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    Odrv12 I__2213 (
            .O(N__21266),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ));
    InMux I__2212 (
            .O(N__21255),
            .I(N__21252));
    LocalMux I__2211 (
            .O(N__21252),
            .I(N__21248));
    InMux I__2210 (
            .O(N__21251),
            .I(N__21245));
    Span4Mux_v I__2209 (
            .O(N__21248),
            .I(N__21240));
    LocalMux I__2208 (
            .O(N__21245),
            .I(N__21240));
    Span4Mux_v I__2207 (
            .O(N__21240),
            .I(N__21237));
    Span4Mux_v I__2206 (
            .O(N__21237),
            .I(N__21234));
    Odrv4 I__2205 (
            .O(N__21234),
            .I(\pwm_generator_inst.un3_threshold_acc ));
    InMux I__2204 (
            .O(N__21231),
            .I(N__21228));
    LocalMux I__2203 (
            .O(N__21228),
            .I(N__21225));
    Odrv4 I__2202 (
            .O(N__21225),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_1 ));
    InMux I__2201 (
            .O(N__21222),
            .I(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ));
    CascadeMux I__2200 (
            .O(N__21219),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    CascadeMux I__2199 (
            .O(N__21216),
            .I(\pwm_generator_inst.un1_counterlto9_2_cascade_ ));
    InMux I__2198 (
            .O(N__21213),
            .I(N__21210));
    LocalMux I__2197 (
            .O(N__21210),
            .I(\pwm_generator_inst.un1_counterlt9 ));
    CascadeMux I__2196 (
            .O(N__21207),
            .I(N__21204));
    InMux I__2195 (
            .O(N__21204),
            .I(N__21201));
    LocalMux I__2194 (
            .O(N__21201),
            .I(N__21198));
    Span4Mux_v I__2193 (
            .O(N__21198),
            .I(N__21194));
    InMux I__2192 (
            .O(N__21197),
            .I(N__21191));
    Odrv4 I__2191 (
            .O(N__21194),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    LocalMux I__2190 (
            .O(N__21191),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ));
    InMux I__2189 (
            .O(N__21186),
            .I(N__21183));
    LocalMux I__2188 (
            .O(N__21183),
            .I(N__21180));
    Span4Mux_h I__2187 (
            .O(N__21180),
            .I(N__21177));
    Span4Mux_v I__2186 (
            .O(N__21177),
            .I(N__21174));
    Span4Mux_v I__2185 (
            .O(N__21174),
            .I(N__21171));
    Odrv4 I__2184 (
            .O(N__21171),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__2183 (
            .O(N__21168),
            .I(N__21165));
    LocalMux I__2182 (
            .O(N__21165),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ));
    InMux I__2181 (
            .O(N__21162),
            .I(N__21159));
    LocalMux I__2180 (
            .O(N__21159),
            .I(N__21156));
    Span4Mux_h I__2179 (
            .O(N__21156),
            .I(N__21153));
    Sp12to4 I__2178 (
            .O(N__21153),
            .I(N__21150));
    Odrv12 I__2177 (
            .O(N__21150),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__2176 (
            .O(N__21147),
            .I(N__21144));
    LocalMux I__2175 (
            .O(N__21144),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ));
    InMux I__2174 (
            .O(N__21141),
            .I(N__21138));
    LocalMux I__2173 (
            .O(N__21138),
            .I(N__21135));
    Span12Mux_h I__2172 (
            .O(N__21135),
            .I(N__21132));
    Odrv12 I__2171 (
            .O(N__21132),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__2170 (
            .O(N__21129),
            .I(N__21126));
    LocalMux I__2169 (
            .O(N__21126),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ));
    InMux I__2168 (
            .O(N__21123),
            .I(N__21120));
    LocalMux I__2167 (
            .O(N__21120),
            .I(N__21117));
    Span4Mux_h I__2166 (
            .O(N__21117),
            .I(N__21114));
    Sp12to4 I__2165 (
            .O(N__21114),
            .I(N__21111));
    Odrv12 I__2164 (
            .O(N__21111),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__2163 (
            .O(N__21108),
            .I(N__21105));
    LocalMux I__2162 (
            .O(N__21105),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ));
    InMux I__2161 (
            .O(N__21102),
            .I(N__21099));
    LocalMux I__2160 (
            .O(N__21099),
            .I(\pwm_generator_inst.thresholdZ0Z_3 ));
    CascadeMux I__2159 (
            .O(N__21096),
            .I(N__21093));
    InMux I__2158 (
            .O(N__21093),
            .I(N__21090));
    LocalMux I__2157 (
            .O(N__21090),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__2156 (
            .O(N__21087),
            .I(N__21084));
    LocalMux I__2155 (
            .O(N__21084),
            .I(N__21081));
    Odrv4 I__2154 (
            .O(N__21081),
            .I(\pwm_generator_inst.thresholdZ0Z_4 ));
    CascadeMux I__2153 (
            .O(N__21078),
            .I(N__21075));
    InMux I__2152 (
            .O(N__21075),
            .I(N__21072));
    LocalMux I__2151 (
            .O(N__21072),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__2150 (
            .O(N__21069),
            .I(N__21066));
    InMux I__2149 (
            .O(N__21066),
            .I(N__21063));
    LocalMux I__2148 (
            .O(N__21063),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__2147 (
            .O(N__21060),
            .I(N__21057));
    InMux I__2146 (
            .O(N__21057),
            .I(N__21054));
    LocalMux I__2145 (
            .O(N__21054),
            .I(\pwm_generator_inst.thresholdZ0Z_6 ));
    InMux I__2144 (
            .O(N__21051),
            .I(N__21048));
    LocalMux I__2143 (
            .O(N__21048),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__2142 (
            .O(N__21045),
            .I(N__21042));
    LocalMux I__2141 (
            .O(N__21042),
            .I(N__21039));
    Odrv4 I__2140 (
            .O(N__21039),
            .I(\pwm_generator_inst.thresholdZ0Z_7 ));
    CascadeMux I__2139 (
            .O(N__21036),
            .I(N__21033));
    InMux I__2138 (
            .O(N__21033),
            .I(N__21030));
    LocalMux I__2137 (
            .O(N__21030),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2136 (
            .O(N__21027),
            .I(N__21024));
    InMux I__2135 (
            .O(N__21024),
            .I(N__21021));
    LocalMux I__2134 (
            .O(N__21021),
            .I(\pwm_generator_inst.counter_i_8 ));
    InMux I__2133 (
            .O(N__21018),
            .I(N__21015));
    LocalMux I__2132 (
            .O(N__21015),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2131 (
            .O(N__21012),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2130 (
            .O(N__21009),
            .I(N__21006));
    LocalMux I__2129 (
            .O(N__21006),
            .I(N__21003));
    Span4Mux_s1_v I__2128 (
            .O(N__21003),
            .I(N__21000));
    Sp12to4 I__2127 (
            .O(N__21000),
            .I(N__20997));
    Span12Mux_s10_h I__2126 (
            .O(N__20997),
            .I(N__20994));
    Span12Mux_h I__2125 (
            .O(N__20994),
            .I(N__20991));
    Odrv12 I__2124 (
            .O(N__20991),
            .I(pwm_output_c));
    CascadeMux I__2123 (
            .O(N__20988),
            .I(N__20985));
    InMux I__2122 (
            .O(N__20985),
            .I(N__20982));
    LocalMux I__2121 (
            .O(N__20982),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ));
    InMux I__2120 (
            .O(N__20979),
            .I(N__20972));
    InMux I__2119 (
            .O(N__20978),
            .I(N__20972));
    CascadeMux I__2118 (
            .O(N__20977),
            .I(N__20969));
    LocalMux I__2117 (
            .O(N__20972),
            .I(N__20963));
    InMux I__2116 (
            .O(N__20969),
            .I(N__20960));
    InMux I__2115 (
            .O(N__20968),
            .I(N__20953));
    InMux I__2114 (
            .O(N__20967),
            .I(N__20953));
    InMux I__2113 (
            .O(N__20966),
            .I(N__20953));
    Span4Mux_v I__2112 (
            .O(N__20963),
            .I(N__20947));
    LocalMux I__2111 (
            .O(N__20960),
            .I(N__20947));
    LocalMux I__2110 (
            .O(N__20953),
            .I(N__20944));
    InMux I__2109 (
            .O(N__20952),
            .I(N__20941));
    Span4Mux_v I__2108 (
            .O(N__20947),
            .I(N__20938));
    Span4Mux_s3_h I__2107 (
            .O(N__20944),
            .I(N__20935));
    LocalMux I__2106 (
            .O(N__20941),
            .I(N__20932));
    Odrv4 I__2105 (
            .O(N__20938),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2104 (
            .O(N__20935),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2103 (
            .O(N__20932),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2102 (
            .O(N__20925),
            .I(N__20922));
    LocalMux I__2101 (
            .O(N__20922),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_1 ));
    InMux I__2100 (
            .O(N__20919),
            .I(N__20916));
    LocalMux I__2099 (
            .O(N__20916),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_3 ));
    InMux I__2098 (
            .O(N__20913),
            .I(N__20910));
    LocalMux I__2097 (
            .O(N__20910),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_2 ));
    CascadeMux I__2096 (
            .O(N__20907),
            .I(N__20904));
    InMux I__2095 (
            .O(N__20904),
            .I(N__20901));
    LocalMux I__2094 (
            .O(N__20901),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__2093 (
            .O(N__20898),
            .I(N__20895));
    LocalMux I__2092 (
            .O(N__20895),
            .I(\pwm_generator_inst.thresholdZ0Z_1 ));
    CascadeMux I__2091 (
            .O(N__20892),
            .I(N__20889));
    InMux I__2090 (
            .O(N__20889),
            .I(N__20886));
    LocalMux I__2089 (
            .O(N__20886),
            .I(\pwm_generator_inst.counter_i_1 ));
    InMux I__2088 (
            .O(N__20883),
            .I(N__20880));
    LocalMux I__2087 (
            .O(N__20880),
            .I(N__20877));
    Odrv4 I__2086 (
            .O(N__20877),
            .I(\pwm_generator_inst.thresholdZ0Z_2 ));
    CascadeMux I__2085 (
            .O(N__20874),
            .I(N__20871));
    InMux I__2084 (
            .O(N__20871),
            .I(N__20868));
    LocalMux I__2083 (
            .O(N__20868),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__2082 (
            .O(N__20865),
            .I(N__20862));
    LocalMux I__2081 (
            .O(N__20862),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_3 ));
    InMux I__2080 (
            .O(N__20859),
            .I(N__20856));
    LocalMux I__2079 (
            .O(N__20856),
            .I(N__20853));
    Odrv12 I__2078 (
            .O(N__20853),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ));
    InMux I__2077 (
            .O(N__20850),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_2 ));
    InMux I__2076 (
            .O(N__20847),
            .I(N__20844));
    LocalMux I__2075 (
            .O(N__20844),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_4 ));
    InMux I__2074 (
            .O(N__20841),
            .I(N__20838));
    LocalMux I__2073 (
            .O(N__20838),
            .I(N__20835));
    Odrv12 I__2072 (
            .O(N__20835),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ));
    InMux I__2071 (
            .O(N__20832),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_3 ));
    InMux I__2070 (
            .O(N__20829),
            .I(N__20826));
    LocalMux I__2069 (
            .O(N__20826),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_5 ));
    InMux I__2068 (
            .O(N__20823),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_4 ));
    InMux I__2067 (
            .O(N__20820),
            .I(N__20817));
    LocalMux I__2066 (
            .O(N__20817),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_6 ));
    CascadeMux I__2065 (
            .O(N__20814),
            .I(N__20811));
    InMux I__2064 (
            .O(N__20811),
            .I(N__20808));
    LocalMux I__2063 (
            .O(N__20808),
            .I(N__20805));
    Span4Mux_v I__2062 (
            .O(N__20805),
            .I(N__20802));
    Odrv4 I__2061 (
            .O(N__20802),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ));
    InMux I__2060 (
            .O(N__20799),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_5 ));
    InMux I__2059 (
            .O(N__20796),
            .I(N__20793));
    LocalMux I__2058 (
            .O(N__20793),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_7 ));
    InMux I__2057 (
            .O(N__20790),
            .I(N__20787));
    LocalMux I__2056 (
            .O(N__20787),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ));
    InMux I__2055 (
            .O(N__20784),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_6 ));
    InMux I__2054 (
            .O(N__20781),
            .I(bfn_2_19_0_));
    InMux I__2053 (
            .O(N__20778),
            .I(N__20775));
    LocalMux I__2052 (
            .O(N__20775),
            .I(N__20772));
    Odrv12 I__2051 (
            .O(N__20772),
            .I(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ));
    InMux I__2050 (
            .O(N__20769),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_8 ));
    CascadeMux I__2049 (
            .O(N__20766),
            .I(N__20763));
    InMux I__2048 (
            .O(N__20763),
            .I(N__20760));
    LocalMux I__2047 (
            .O(N__20760),
            .I(N__20756));
    InMux I__2046 (
            .O(N__20759),
            .I(N__20753));
    Span4Mux_v I__2045 (
            .O(N__20756),
            .I(N__20748));
    LocalMux I__2044 (
            .O(N__20753),
            .I(N__20748));
    Odrv4 I__2043 (
            .O(N__20748),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ));
    InMux I__2042 (
            .O(N__20745),
            .I(N__20742));
    LocalMux I__2041 (
            .O(N__20742),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_8 ));
    CascadeMux I__2040 (
            .O(N__20739),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ));
    InMux I__2039 (
            .O(N__20736),
            .I(N__20730));
    InMux I__2038 (
            .O(N__20735),
            .I(N__20730));
    LocalMux I__2037 (
            .O(N__20730),
            .I(N__20727));
    Odrv4 I__2036 (
            .O(N__20727),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ));
    InMux I__2035 (
            .O(N__20724),
            .I(N__20718));
    InMux I__2034 (
            .O(N__20723),
            .I(N__20718));
    LocalMux I__2033 (
            .O(N__20718),
            .I(N__20715));
    Odrv4 I__2032 (
            .O(N__20715),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ));
    CascadeMux I__2031 (
            .O(N__20712),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ));
    InMux I__2030 (
            .O(N__20709),
            .I(N__20703));
    InMux I__2029 (
            .O(N__20708),
            .I(N__20703));
    LocalMux I__2028 (
            .O(N__20703),
            .I(N__20700));
    Odrv4 I__2027 (
            .O(N__20700),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ));
    CascadeMux I__2026 (
            .O(N__20697),
            .I(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ));
    CascadeMux I__2025 (
            .O(N__20694),
            .I(N__20691));
    InMux I__2024 (
            .O(N__20691),
            .I(N__20687));
    InMux I__2023 (
            .O(N__20690),
            .I(N__20684));
    LocalMux I__2022 (
            .O(N__20687),
            .I(N__20679));
    LocalMux I__2021 (
            .O(N__20684),
            .I(N__20679));
    Odrv4 I__2020 (
            .O(N__20679),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ));
    InMux I__2019 (
            .O(N__20676),
            .I(N__20673));
    LocalMux I__2018 (
            .O(N__20673),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_0 ));
    CascadeMux I__2017 (
            .O(N__20670),
            .I(N__20667));
    InMux I__2016 (
            .O(N__20667),
            .I(N__20664));
    LocalMux I__2015 (
            .O(N__20664),
            .I(N__20661));
    Odrv12 I__2014 (
            .O(N__20661),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ));
    InMux I__2013 (
            .O(N__20658),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_0 ));
    InMux I__2012 (
            .O(N__20655),
            .I(N__20652));
    LocalMux I__2011 (
            .O(N__20652),
            .I(\pwm_generator_inst.un19_threshold_acc_axb_2 ));
    CascadeMux I__2010 (
            .O(N__20649),
            .I(N__20646));
    InMux I__2009 (
            .O(N__20646),
            .I(N__20643));
    LocalMux I__2008 (
            .O(N__20643),
            .I(N__20640));
    Odrv12 I__2007 (
            .O(N__20640),
            .I(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ));
    InMux I__2006 (
            .O(N__20637),
            .I(\pwm_generator_inst.un19_threshold_acc_cry_1 ));
    InMux I__2005 (
            .O(N__20634),
            .I(N__20631));
    LocalMux I__2004 (
            .O(N__20631),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ));
    InMux I__2003 (
            .O(N__20628),
            .I(N__20625));
    LocalMux I__2002 (
            .O(N__20625),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ));
    InMux I__2001 (
            .O(N__20622),
            .I(N__20619));
    LocalMux I__2000 (
            .O(N__20619),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ));
    InMux I__1999 (
            .O(N__20616),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19 ));
    InMux I__1998 (
            .O(N__20613),
            .I(N__20610));
    LocalMux I__1997 (
            .O(N__20610),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ));
    CascadeMux I__1996 (
            .O(N__20607),
            .I(N__20604));
    InMux I__1995 (
            .O(N__20604),
            .I(N__20601));
    LocalMux I__1994 (
            .O(N__20601),
            .I(N__20597));
    InMux I__1993 (
            .O(N__20600),
            .I(N__20594));
    Span4Mux_v I__1992 (
            .O(N__20597),
            .I(N__20589));
    LocalMux I__1991 (
            .O(N__20594),
            .I(N__20589));
    Odrv4 I__1990 (
            .O(N__20589),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ));
    InMux I__1989 (
            .O(N__20586),
            .I(N__20583));
    LocalMux I__1988 (
            .O(N__20583),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ));
    InMux I__1987 (
            .O(N__20580),
            .I(bfn_2_15_0_));
    InMux I__1986 (
            .O(N__20577),
            .I(N__20574));
    LocalMux I__1985 (
            .O(N__20574),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ));
    InMux I__1984 (
            .O(N__20571),
            .I(N__20568));
    LocalMux I__1983 (
            .O(N__20568),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ));
    InMux I__1982 (
            .O(N__20565),
            .I(N__20562));
    LocalMux I__1981 (
            .O(N__20562),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ));
    InMux I__1980 (
            .O(N__20559),
            .I(N__20556));
    LocalMux I__1979 (
            .O(N__20556),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ));
    InMux I__1978 (
            .O(N__20553),
            .I(N__20550));
    LocalMux I__1977 (
            .O(N__20550),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ));
    InMux I__1976 (
            .O(N__20547),
            .I(N__20544));
    LocalMux I__1975 (
            .O(N__20544),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ));
    InMux I__1974 (
            .O(N__20541),
            .I(N__20538));
    LocalMux I__1973 (
            .O(N__20538),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ));
    InMux I__1972 (
            .O(N__20535),
            .I(N__20532));
    LocalMux I__1971 (
            .O(N__20532),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ));
    InMux I__1970 (
            .O(N__20529),
            .I(N__20526));
    LocalMux I__1969 (
            .O(N__20526),
            .I(N__20523));
    Span4Mux_v I__1968 (
            .O(N__20523),
            .I(N__20520));
    Span4Mux_v I__1967 (
            .O(N__20520),
            .I(N__20517));
    Odrv4 I__1966 (
            .O(N__20517),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1965 (
            .O(N__20514),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_0 ));
    InMux I__1964 (
            .O(N__20511),
            .I(N__20508));
    LocalMux I__1963 (
            .O(N__20508),
            .I(N__20505));
    Span4Mux_v I__1962 (
            .O(N__20505),
            .I(N__20502));
    Span4Mux_v I__1961 (
            .O(N__20502),
            .I(N__20499));
    Odrv4 I__1960 (
            .O(N__20499),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1959 (
            .O(N__20496),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_1 ));
    InMux I__1958 (
            .O(N__20493),
            .I(N__20490));
    LocalMux I__1957 (
            .O(N__20490),
            .I(N__20487));
    Span12Mux_v I__1956 (
            .O(N__20487),
            .I(N__20484));
    Odrv12 I__1955 (
            .O(N__20484),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1954 (
            .O(N__20481),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_2 ));
    InMux I__1953 (
            .O(N__20478),
            .I(N__20475));
    LocalMux I__1952 (
            .O(N__20475),
            .I(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ));
    InMux I__1951 (
            .O(N__20472),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_3 ));
    CascadeMux I__1950 (
            .O(N__20469),
            .I(N__20466));
    InMux I__1949 (
            .O(N__20466),
            .I(N__20463));
    LocalMux I__1948 (
            .O(N__20463),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ));
    InMux I__1947 (
            .O(N__20460),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_4 ));
    CascadeMux I__1946 (
            .O(N__20457),
            .I(N__20454));
    InMux I__1945 (
            .O(N__20454),
            .I(N__20451));
    LocalMux I__1944 (
            .O(N__20451),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ));
    InMux I__1943 (
            .O(N__20448),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_5 ));
    CascadeMux I__1942 (
            .O(N__20445),
            .I(N__20442));
    InMux I__1941 (
            .O(N__20442),
            .I(N__20439));
    LocalMux I__1940 (
            .O(N__20439),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ));
    InMux I__1939 (
            .O(N__20436),
            .I(\pwm_generator_inst.un3_threshold_acc_cry_6 ));
    CascadeMux I__1938 (
            .O(N__20433),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    CascadeMux I__1937 (
            .O(N__20430),
            .I(N__20426));
    CascadeMux I__1936 (
            .O(N__20429),
            .I(N__20423));
    InMux I__1935 (
            .O(N__20426),
            .I(N__20420));
    InMux I__1934 (
            .O(N__20423),
            .I(N__20417));
    LocalMux I__1933 (
            .O(N__20420),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__1932 (
            .O(N__20417),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__1931 (
            .O(N__20412),
            .I(\current_shift_inst.PI_CTRL.N_31_cascade_ ));
    InMux I__1930 (
            .O(N__20409),
            .I(N__20405));
    InMux I__1929 (
            .O(N__20408),
            .I(N__20402));
    LocalMux I__1928 (
            .O(N__20405),
            .I(N__20397));
    LocalMux I__1927 (
            .O(N__20402),
            .I(N__20397));
    Odrv4 I__1926 (
            .O(N__20397),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    InMux I__1925 (
            .O(N__20394),
            .I(N__20391));
    LocalMux I__1924 (
            .O(N__20391),
            .I(N__20388));
    Span12Mux_v I__1923 (
            .O(N__20388),
            .I(N__20385));
    Odrv12 I__1922 (
            .O(N__20385),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_7 ));
    InMux I__1921 (
            .O(N__20382),
            .I(N__20379));
    LocalMux I__1920 (
            .O(N__20379),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_6 ));
    InMux I__1919 (
            .O(N__20376),
            .I(N__20373));
    LocalMux I__1918 (
            .O(N__20373),
            .I(\pwm_generator_inst.threshold_ACCZ0Z_4 ));
    InMux I__1917 (
            .O(N__20370),
            .I(N__20363));
    InMux I__1916 (
            .O(N__20369),
            .I(N__20363));
    InMux I__1915 (
            .O(N__20368),
            .I(N__20360));
    LocalMux I__1914 (
            .O(N__20363),
            .I(pwm_duty_input_8));
    LocalMux I__1913 (
            .O(N__20360),
            .I(pwm_duty_input_8));
    InMux I__1912 (
            .O(N__20355),
            .I(N__20348));
    InMux I__1911 (
            .O(N__20354),
            .I(N__20348));
    InMux I__1910 (
            .O(N__20353),
            .I(N__20345));
    LocalMux I__1909 (
            .O(N__20348),
            .I(pwm_duty_input_9));
    LocalMux I__1908 (
            .O(N__20345),
            .I(pwm_duty_input_9));
    CascadeMux I__1907 (
            .O(N__20340),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__1906 (
            .O(N__20337),
            .I(N__20334));
    LocalMux I__1905 (
            .O(N__20334),
            .I(N__20329));
    InMux I__1904 (
            .O(N__20333),
            .I(N__20324));
    InMux I__1903 (
            .O(N__20332),
            .I(N__20324));
    Span4Mux_s1_h I__1902 (
            .O(N__20329),
            .I(N__20321));
    LocalMux I__1901 (
            .O(N__20324),
            .I(pwm_duty_input_6));
    Odrv4 I__1900 (
            .O(N__20321),
            .I(pwm_duty_input_6));
    InMux I__1899 (
            .O(N__20316),
            .I(N__20313));
    LocalMux I__1898 (
            .O(N__20313),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__1897 (
            .O(N__20310),
            .I(\current_shift_inst.PI_CTRL.N_27_cascade_ ));
    CascadeMux I__1896 (
            .O(N__20307),
            .I(N__20301));
    CascadeMux I__1895 (
            .O(N__20306),
            .I(N__20298));
    CascadeMux I__1894 (
            .O(N__20305),
            .I(N__20295));
    CascadeMux I__1893 (
            .O(N__20304),
            .I(N__20292));
    InMux I__1892 (
            .O(N__20301),
            .I(N__20287));
    InMux I__1891 (
            .O(N__20298),
            .I(N__20287));
    InMux I__1890 (
            .O(N__20295),
            .I(N__20283));
    InMux I__1889 (
            .O(N__20292),
            .I(N__20280));
    LocalMux I__1888 (
            .O(N__20287),
            .I(N__20277));
    InMux I__1887 (
            .O(N__20286),
            .I(N__20274));
    LocalMux I__1886 (
            .O(N__20283),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    LocalMux I__1885 (
            .O(N__20280),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    Odrv4 I__1884 (
            .O(N__20277),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    LocalMux I__1883 (
            .O(N__20274),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    CascadeMux I__1882 (
            .O(N__20265),
            .I(N__20262));
    InMux I__1881 (
            .O(N__20262),
            .I(N__20258));
    InMux I__1880 (
            .O(N__20261),
            .I(N__20255));
    LocalMux I__1879 (
            .O(N__20258),
            .I(N__20251));
    LocalMux I__1878 (
            .O(N__20255),
            .I(N__20248));
    InMux I__1877 (
            .O(N__20254),
            .I(N__20245));
    Span4Mux_h I__1876 (
            .O(N__20251),
            .I(N__20240));
    Span4Mux_s1_h I__1875 (
            .O(N__20248),
            .I(N__20240));
    LocalMux I__1874 (
            .O(N__20245),
            .I(pwm_duty_input_5));
    Odrv4 I__1873 (
            .O(N__20240),
            .I(pwm_duty_input_5));
    InMux I__1872 (
            .O(N__20235),
            .I(N__20232));
    LocalMux I__1871 (
            .O(N__20232),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    InMux I__1870 (
            .O(N__20229),
            .I(N__20226));
    LocalMux I__1869 (
            .O(N__20226),
            .I(N__20223));
    Odrv4 I__1868 (
            .O(N__20223),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    InMux I__1867 (
            .O(N__20220),
            .I(N__20213));
    InMux I__1866 (
            .O(N__20219),
            .I(N__20213));
    InMux I__1865 (
            .O(N__20218),
            .I(N__20210));
    LocalMux I__1864 (
            .O(N__20213),
            .I(pwm_duty_input_4));
    LocalMux I__1863 (
            .O(N__20210),
            .I(pwm_duty_input_4));
    CascadeMux I__1862 (
            .O(N__20205),
            .I(N__20201));
    InMux I__1861 (
            .O(N__20204),
            .I(N__20197));
    InMux I__1860 (
            .O(N__20201),
            .I(N__20192));
    InMux I__1859 (
            .O(N__20200),
            .I(N__20192));
    LocalMux I__1858 (
            .O(N__20197),
            .I(N__20189));
    LocalMux I__1857 (
            .O(N__20192),
            .I(pwm_duty_input_3));
    Odrv4 I__1856 (
            .O(N__20189),
            .I(pwm_duty_input_3));
    InMux I__1855 (
            .O(N__20184),
            .I(N__20181));
    LocalMux I__1854 (
            .O(N__20181),
            .I(N__20178));
    Odrv4 I__1853 (
            .O(N__20178),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__1852 (
            .O(N__20175),
            .I(N__20169));
    InMux I__1851 (
            .O(N__20174),
            .I(N__20169));
    LocalMux I__1850 (
            .O(N__20169),
            .I(N__20165));
    InMux I__1849 (
            .O(N__20168),
            .I(N__20162));
    Odrv4 I__1848 (
            .O(N__20165),
            .I(\current_shift_inst.PI_CTRL.N_154 ));
    LocalMux I__1847 (
            .O(N__20162),
            .I(\current_shift_inst.PI_CTRL.N_154 ));
    InMux I__1846 (
            .O(N__20157),
            .I(N__20154));
    LocalMux I__1845 (
            .O(N__20154),
            .I(\current_shift_inst.PI_CTRL.N_155 ));
    InMux I__1844 (
            .O(N__20151),
            .I(bfn_1_16_0_));
    InMux I__1843 (
            .O(N__20148),
            .I(N__20145));
    LocalMux I__1842 (
            .O(N__20145),
            .I(un7_start_stop_0_a2));
    InMux I__1841 (
            .O(N__20142),
            .I(N__20139));
    LocalMux I__1840 (
            .O(N__20139),
            .I(N_38_i_i));
    InMux I__1839 (
            .O(N__20136),
            .I(N__20132));
    InMux I__1838 (
            .O(N__20135),
            .I(N__20129));
    LocalMux I__1837 (
            .O(N__20132),
            .I(N__20126));
    LocalMux I__1836 (
            .O(N__20129),
            .I(pwm_duty_input_0));
    Odrv4 I__1835 (
            .O(N__20126),
            .I(pwm_duty_input_0));
    InMux I__1834 (
            .O(N__20121),
            .I(N__20117));
    InMux I__1833 (
            .O(N__20120),
            .I(N__20114));
    LocalMux I__1832 (
            .O(N__20117),
            .I(N__20111));
    LocalMux I__1831 (
            .O(N__20114),
            .I(pwm_duty_input_1));
    Odrv4 I__1830 (
            .O(N__20111),
            .I(pwm_duty_input_1));
    InMux I__1829 (
            .O(N__20106),
            .I(N__20102));
    InMux I__1828 (
            .O(N__20105),
            .I(N__20099));
    LocalMux I__1827 (
            .O(N__20102),
            .I(pwm_duty_input_2));
    LocalMux I__1826 (
            .O(N__20099),
            .I(pwm_duty_input_2));
    InMux I__1825 (
            .O(N__20094),
            .I(N__20087));
    InMux I__1824 (
            .O(N__20093),
            .I(N__20087));
    InMux I__1823 (
            .O(N__20092),
            .I(N__20084));
    LocalMux I__1822 (
            .O(N__20087),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    LocalMux I__1821 (
            .O(N__20084),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1820 (
            .O(N__20079),
            .I(N__20075));
    CascadeMux I__1819 (
            .O(N__20078),
            .I(N__20072));
    LocalMux I__1818 (
            .O(N__20075),
            .I(N__20068));
    InMux I__1817 (
            .O(N__20072),
            .I(N__20063));
    InMux I__1816 (
            .O(N__20071),
            .I(N__20063));
    Span4Mux_s2_h I__1815 (
            .O(N__20068),
            .I(N__20060));
    LocalMux I__1814 (
            .O(N__20063),
            .I(pwm_duty_input_7));
    Odrv4 I__1813 (
            .O(N__20060),
            .I(pwm_duty_input_7));
    InMux I__1812 (
            .O(N__20055),
            .I(N__20052));
    LocalMux I__1811 (
            .O(N__20052),
            .I(N__20049));
    Span4Mux_v I__1810 (
            .O(N__20049),
            .I(N__20046));
    Odrv4 I__1809 (
            .O(N__20046),
            .I(\pwm_generator_inst.un2_threshold_acc_2_8 ));
    CascadeMux I__1808 (
            .O(N__20043),
            .I(N__20040));
    InMux I__1807 (
            .O(N__20040),
            .I(N__20037));
    LocalMux I__1806 (
            .O(N__20037),
            .I(N__20034));
    Span4Mux_v I__1805 (
            .O(N__20034),
            .I(N__20031));
    Span4Mux_v I__1804 (
            .O(N__20031),
            .I(N__20028));
    Odrv4 I__1803 (
            .O(N__20028),
            .I(\pwm_generator_inst.un2_threshold_acc_1_23 ));
    InMux I__1802 (
            .O(N__20025),
            .I(bfn_1_15_0_));
    InMux I__1801 (
            .O(N__20022),
            .I(N__20019));
    LocalMux I__1800 (
            .O(N__20019),
            .I(N__20016));
    Span4Mux_v I__1799 (
            .O(N__20016),
            .I(N__20013));
    Odrv4 I__1798 (
            .O(N__20013),
            .I(\pwm_generator_inst.un2_threshold_acc_2_9 ));
    CascadeMux I__1797 (
            .O(N__20010),
            .I(N__20007));
    InMux I__1796 (
            .O(N__20007),
            .I(N__20004));
    LocalMux I__1795 (
            .O(N__20004),
            .I(N__20001));
    Span4Mux_v I__1794 (
            .O(N__20001),
            .I(N__19998));
    Span4Mux_v I__1793 (
            .O(N__19998),
            .I(N__19995));
    Odrv4 I__1792 (
            .O(N__19995),
            .I(\pwm_generator_inst.un2_threshold_acc_1_24 ));
    InMux I__1791 (
            .O(N__19992),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ));
    InMux I__1790 (
            .O(N__19989),
            .I(N__19986));
    LocalMux I__1789 (
            .O(N__19986),
            .I(N__19983));
    Span4Mux_v I__1788 (
            .O(N__19983),
            .I(N__19980));
    Odrv4 I__1787 (
            .O(N__19980),
            .I(\pwm_generator_inst.un2_threshold_acc_2_10 ));
    InMux I__1786 (
            .O(N__19977),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ));
    CascadeMux I__1785 (
            .O(N__19974),
            .I(N__19971));
    InMux I__1784 (
            .O(N__19971),
            .I(N__19968));
    LocalMux I__1783 (
            .O(N__19968),
            .I(N__19965));
    Span4Mux_v I__1782 (
            .O(N__19965),
            .I(N__19962));
    Odrv4 I__1781 (
            .O(N__19962),
            .I(\pwm_generator_inst.un2_threshold_acc_2_11 ));
    InMux I__1780 (
            .O(N__19959),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ));
    InMux I__1779 (
            .O(N__19956),
            .I(N__19953));
    LocalMux I__1778 (
            .O(N__19953),
            .I(N__19950));
    Span4Mux_v I__1777 (
            .O(N__19950),
            .I(N__19947));
    Odrv4 I__1776 (
            .O(N__19947),
            .I(\pwm_generator_inst.un2_threshold_acc_2_12 ));
    InMux I__1775 (
            .O(N__19944),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ));
    CascadeMux I__1774 (
            .O(N__19941),
            .I(N__19938));
    InMux I__1773 (
            .O(N__19938),
            .I(N__19935));
    LocalMux I__1772 (
            .O(N__19935),
            .I(N__19932));
    Span4Mux_v I__1771 (
            .O(N__19932),
            .I(N__19929));
    Odrv4 I__1770 (
            .O(N__19929),
            .I(\pwm_generator_inst.un2_threshold_acc_2_13 ));
    InMux I__1769 (
            .O(N__19926),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ));
    InMux I__1768 (
            .O(N__19923),
            .I(N__19920));
    LocalMux I__1767 (
            .O(N__19920),
            .I(N__19917));
    Span4Mux_v I__1766 (
            .O(N__19917),
            .I(N__19914));
    Odrv4 I__1765 (
            .O(N__19914),
            .I(\pwm_generator_inst.un2_threshold_acc_2_14 ));
    InMux I__1764 (
            .O(N__19911),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ));
    CascadeMux I__1763 (
            .O(N__19908),
            .I(N__19902));
    CascadeMux I__1762 (
            .O(N__19907),
            .I(N__19898));
    CascadeMux I__1761 (
            .O(N__19906),
            .I(N__19894));
    InMux I__1760 (
            .O(N__19905),
            .I(N__19879));
    InMux I__1759 (
            .O(N__19902),
            .I(N__19879));
    InMux I__1758 (
            .O(N__19901),
            .I(N__19879));
    InMux I__1757 (
            .O(N__19898),
            .I(N__19879));
    InMux I__1756 (
            .O(N__19897),
            .I(N__19879));
    InMux I__1755 (
            .O(N__19894),
            .I(N__19879));
    InMux I__1754 (
            .O(N__19893),
            .I(N__19876));
    InMux I__1753 (
            .O(N__19892),
            .I(N__19873));
    LocalMux I__1752 (
            .O(N__19879),
            .I(N__19870));
    LocalMux I__1751 (
            .O(N__19876),
            .I(N__19867));
    LocalMux I__1750 (
            .O(N__19873),
            .I(N__19862));
    Span4Mux_v I__1749 (
            .O(N__19870),
            .I(N__19862));
    Span4Mux_v I__1748 (
            .O(N__19867),
            .I(N__19857));
    Span4Mux_v I__1747 (
            .O(N__19862),
            .I(N__19857));
    Odrv4 I__1746 (
            .O(N__19857),
            .I(\pwm_generator_inst.un2_threshold_acc_1_25 ));
    CascadeMux I__1745 (
            .O(N__19854),
            .I(N__19851));
    InMux I__1744 (
            .O(N__19851),
            .I(N__19848));
    LocalMux I__1743 (
            .O(N__19848),
            .I(N__19845));
    Odrv12 I__1742 (
            .O(N__19845),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ));
    InMux I__1741 (
            .O(N__19842),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ));
    InMux I__1740 (
            .O(N__19839),
            .I(N__19836));
    LocalMux I__1739 (
            .O(N__19836),
            .I(N__19833));
    Odrv12 I__1738 (
            .O(N__19833),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ));
    InMux I__1737 (
            .O(N__19830),
            .I(N__19827));
    LocalMux I__1736 (
            .O(N__19827),
            .I(N__19824));
    Span4Mux_v I__1735 (
            .O(N__19824),
            .I(N__19821));
    Odrv4 I__1734 (
            .O(N__19821),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1 ));
    CascadeMux I__1733 (
            .O(N__19818),
            .I(N__19815));
    InMux I__1732 (
            .O(N__19815),
            .I(N__19812));
    LocalMux I__1731 (
            .O(N__19812),
            .I(N__19809));
    Span4Mux_v I__1730 (
            .O(N__19809),
            .I(N__19806));
    Span4Mux_v I__1729 (
            .O(N__19806),
            .I(N__19803));
    Odrv4 I__1728 (
            .O(N__19803),
            .I(\pwm_generator_inst.un2_threshold_acc_1_16 ));
    InMux I__1727 (
            .O(N__19800),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ));
    InMux I__1726 (
            .O(N__19797),
            .I(N__19794));
    LocalMux I__1725 (
            .O(N__19794),
            .I(N__19791));
    Span4Mux_v I__1724 (
            .O(N__19791),
            .I(N__19788));
    Odrv4 I__1723 (
            .O(N__19788),
            .I(\pwm_generator_inst.un2_threshold_acc_2_2 ));
    CascadeMux I__1722 (
            .O(N__19785),
            .I(N__19782));
    InMux I__1721 (
            .O(N__19782),
            .I(N__19779));
    LocalMux I__1720 (
            .O(N__19779),
            .I(N__19776));
    Span4Mux_v I__1719 (
            .O(N__19776),
            .I(N__19773));
    Span4Mux_v I__1718 (
            .O(N__19773),
            .I(N__19770));
    Odrv4 I__1717 (
            .O(N__19770),
            .I(\pwm_generator_inst.un2_threshold_acc_1_17 ));
    InMux I__1716 (
            .O(N__19767),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ));
    InMux I__1715 (
            .O(N__19764),
            .I(N__19761));
    LocalMux I__1714 (
            .O(N__19761),
            .I(N__19758));
    Span4Mux_v I__1713 (
            .O(N__19758),
            .I(N__19755));
    Odrv4 I__1712 (
            .O(N__19755),
            .I(\pwm_generator_inst.un2_threshold_acc_2_3 ));
    CascadeMux I__1711 (
            .O(N__19752),
            .I(N__19749));
    InMux I__1710 (
            .O(N__19749),
            .I(N__19746));
    LocalMux I__1709 (
            .O(N__19746),
            .I(N__19743));
    Span4Mux_v I__1708 (
            .O(N__19743),
            .I(N__19740));
    Odrv4 I__1707 (
            .O(N__19740),
            .I(\pwm_generator_inst.un2_threshold_acc_1_18 ));
    InMux I__1706 (
            .O(N__19737),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ));
    InMux I__1705 (
            .O(N__19734),
            .I(N__19731));
    LocalMux I__1704 (
            .O(N__19731),
            .I(N__19728));
    Span4Mux_v I__1703 (
            .O(N__19728),
            .I(N__19725));
    Odrv4 I__1702 (
            .O(N__19725),
            .I(\pwm_generator_inst.un2_threshold_acc_2_4 ));
    CascadeMux I__1701 (
            .O(N__19722),
            .I(N__19719));
    InMux I__1700 (
            .O(N__19719),
            .I(N__19716));
    LocalMux I__1699 (
            .O(N__19716),
            .I(N__19713));
    Span4Mux_h I__1698 (
            .O(N__19713),
            .I(N__19710));
    Span4Mux_v I__1697 (
            .O(N__19710),
            .I(N__19707));
    Odrv4 I__1696 (
            .O(N__19707),
            .I(\pwm_generator_inst.un2_threshold_acc_1_19 ));
    InMux I__1695 (
            .O(N__19704),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ));
    InMux I__1694 (
            .O(N__19701),
            .I(N__19698));
    LocalMux I__1693 (
            .O(N__19698),
            .I(N__19695));
    Span4Mux_v I__1692 (
            .O(N__19695),
            .I(N__19692));
    Odrv4 I__1691 (
            .O(N__19692),
            .I(\pwm_generator_inst.un2_threshold_acc_2_5 ));
    CascadeMux I__1690 (
            .O(N__19689),
            .I(N__19686));
    InMux I__1689 (
            .O(N__19686),
            .I(N__19683));
    LocalMux I__1688 (
            .O(N__19683),
            .I(N__19680));
    Span4Mux_v I__1687 (
            .O(N__19680),
            .I(N__19677));
    Odrv4 I__1686 (
            .O(N__19677),
            .I(\pwm_generator_inst.un2_threshold_acc_1_20 ));
    InMux I__1685 (
            .O(N__19674),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ));
    InMux I__1684 (
            .O(N__19671),
            .I(N__19668));
    LocalMux I__1683 (
            .O(N__19668),
            .I(N__19665));
    Span4Mux_v I__1682 (
            .O(N__19665),
            .I(N__19662));
    Odrv4 I__1681 (
            .O(N__19662),
            .I(\pwm_generator_inst.un2_threshold_acc_2_6 ));
    CascadeMux I__1680 (
            .O(N__19659),
            .I(N__19656));
    InMux I__1679 (
            .O(N__19656),
            .I(N__19653));
    LocalMux I__1678 (
            .O(N__19653),
            .I(N__19650));
    Span4Mux_v I__1677 (
            .O(N__19650),
            .I(N__19647));
    Odrv4 I__1676 (
            .O(N__19647),
            .I(\pwm_generator_inst.un2_threshold_acc_1_21 ));
    InMux I__1675 (
            .O(N__19644),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ));
    InMux I__1674 (
            .O(N__19641),
            .I(N__19638));
    LocalMux I__1673 (
            .O(N__19638),
            .I(N__19635));
    Span4Mux_v I__1672 (
            .O(N__19635),
            .I(N__19632));
    Odrv4 I__1671 (
            .O(N__19632),
            .I(\pwm_generator_inst.un2_threshold_acc_2_7 ));
    CascadeMux I__1670 (
            .O(N__19629),
            .I(N__19626));
    InMux I__1669 (
            .O(N__19626),
            .I(N__19623));
    LocalMux I__1668 (
            .O(N__19623),
            .I(N__19620));
    Span4Mux_v I__1667 (
            .O(N__19620),
            .I(N__19617));
    Odrv4 I__1666 (
            .O(N__19617),
            .I(\pwm_generator_inst.un2_threshold_acc_1_22 ));
    InMux I__1665 (
            .O(N__19614),
            .I(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ));
    InMux I__1664 (
            .O(N__19611),
            .I(N__19608));
    LocalMux I__1663 (
            .O(N__19608),
            .I(N__19605));
    Odrv12 I__1662 (
            .O(N__19605),
            .I(\current_shift_inst.PI_CTRL.N_149 ));
    InMux I__1661 (
            .O(N__19602),
            .I(N__19599));
    LocalMux I__1660 (
            .O(N__19599),
            .I(N__19596));
    Odrv4 I__1659 (
            .O(N__19596),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_16 ));
    InMux I__1658 (
            .O(N__19593),
            .I(N__19589));
    InMux I__1657 (
            .O(N__19592),
            .I(N__19586));
    LocalMux I__1656 (
            .O(N__19589),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    LocalMux I__1655 (
            .O(N__19586),
            .I(\pwm_generator_inst.un2_threshold_acc_2_1_15 ));
    InMux I__1654 (
            .O(N__19581),
            .I(N__19578));
    LocalMux I__1653 (
            .O(N__19578),
            .I(N__19575));
    Span4Mux_v I__1652 (
            .O(N__19575),
            .I(N__19572));
    Odrv4 I__1651 (
            .O(N__19572),
            .I(\pwm_generator_inst.un2_threshold_acc_2_0 ));
    CascadeMux I__1650 (
            .O(N__19569),
            .I(N__19566));
    InMux I__1649 (
            .O(N__19566),
            .I(N__19563));
    LocalMux I__1648 (
            .O(N__19563),
            .I(N__19560));
    Span4Mux_v I__1647 (
            .O(N__19560),
            .I(N__19557));
    Span4Mux_v I__1646 (
            .O(N__19557),
            .I(N__19554));
    Odrv4 I__1645 (
            .O(N__19554),
            .I(\pwm_generator_inst.un2_threshold_acc_1_15 ));
    IoInMux I__1644 (
            .O(N__19551),
            .I(N__19548));
    LocalMux I__1643 (
            .O(N__19548),
            .I(N__19545));
    Span4Mux_s3_v I__1642 (
            .O(N__19545),
            .I(N__19542));
    Span4Mux_h I__1641 (
            .O(N__19542),
            .I(N__19539));
    Sp12to4 I__1640 (
            .O(N__19539),
            .I(N__19536));
    Span12Mux_v I__1639 (
            .O(N__19536),
            .I(N__19533));
    Span12Mux_v I__1638 (
            .O(N__19533),
            .I(N__19530));
    Odrv12 I__1637 (
            .O(N__19530),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1636 (
            .O(N__19527),
            .I(N__19524));
    LocalMux I__1635 (
            .O(N__19524),
            .I(N__19521));
    IoSpan4Mux I__1634 (
            .O(N__19521),
            .I(N__19518));
    IoSpan4Mux I__1633 (
            .O(N__19518),
            .I(N__19515));
    Odrv4 I__1632 (
            .O(N__19515),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_8_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_23_0_));
    defparam IN_MUX_bfv_8_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_24_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_8_24_0_));
    defparam IN_MUX_bfv_8_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_25_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_8_25_0_));
    defparam IN_MUX_bfv_8_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_26_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_8_26_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_11_0_));
    defparam IN_MUX_bfv_3_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_12_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_3_12_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_2_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_19_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .carryinitout(bfn_2_19_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_17_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_17_22_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_12_11_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19551),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19527),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__23451),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_393_i_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__35826),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_166_i_g ));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__32016),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_395_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__38270),
            .CLKHFEN(N__38274),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__38283),
            .RGB2PWM(N__20142),
            .RGB1(rgb_g),
            .CURREN(N__38236),
            .RGB2(rgb_b),
            .RGB1PWM(N__20148),
            .RGB0PWM(N__48591),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_1 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_5_1  (
            .in0(N__22203),
            .in1(N__23097),
            .in2(N__22593),
            .in3(N__20979),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49251),
            .ce(),
            .sr(N__48464));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2  (
            .in0(N__20175),
            .in1(N__22737),
            .in2(N__20307),
            .in3(N__20094),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49251),
            .ce(),
            .sr(N__48464));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_6  (
            .in0(N__20174),
            .in1(N__22758),
            .in2(N__20306),
            .in3(N__20093),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49251),
            .ce(),
            .sr(N__48464));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_7 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_5_7  (
            .in0(N__22202),
            .in1(N__23096),
            .in2(N__22632),
            .in3(N__20978),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49251),
            .ce(),
            .sr(N__48464));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_0 .LUT_INIT=16'b1100111111001101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_0  (
            .in0(N__20409),
            .in1(N__22707),
            .in2(N__20304),
            .in3(N__22194),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49250),
            .ce(),
            .sr(N__48470));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_1 .LUT_INIT=16'b1101110001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_6_1  (
            .in0(N__23090),
            .in1(N__22854),
            .in2(N__22201),
            .in3(N__20968),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49250),
            .ce(),
            .sr(N__48470));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2 .LUT_INIT=16'b1011001110110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2  (
            .in0(N__20967),
            .in1(N__23089),
            .in2(N__22923),
            .in3(N__22193),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49250),
            .ce(),
            .sr(N__48470));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_5 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_6_5  (
            .in0(N__20168),
            .in1(N__22722),
            .in2(N__20305),
            .in3(N__20092),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49250),
            .ce(),
            .sr(N__48470));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_6 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_6  (
            .in0(N__20966),
            .in1(N__20316),
            .in2(N__22671),
            .in3(N__19611),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49250),
            .ce(),
            .sr(N__48470));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_7_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_7_0 .LUT_INIT=16'b1010000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_7_0  (
            .in0(N__22886),
            .in1(N__22185),
            .in2(N__20977),
            .in3(N__23088),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49249),
            .ce(),
            .sr(N__48476));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_8_5 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_8_5  (
            .in0(N__23086),
            .in1(N__22664),
            .in2(N__20430),
            .in3(N__22186),
            .lcout(\current_shift_inst.PI_CTRL.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23087),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49247),
            .ce(),
            .sr(N__48497));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_10_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_10_6 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_LC_1_10_6  (
            .in0(N__19593),
            .in1(N__19602),
            .in2(N__21893),
            .in3(N__19892),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofx_LC_1_11_3  (
            .in0(N__19592),
            .in1(N__19893),
            .in2(_gnd_net_),
            .in3(N__21927),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_14_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_axb_4_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__19581),
            .in2(N__19569),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_acc_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_1_s_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__19830),
            .in2(N__19818),
            .in3(N__19800),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_2_s_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__19797),
            .in2(N__19785),
            .in3(N__19767),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_3_s_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__19764),
            .in2(N__19752),
            .in3(N__19737),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_4_s_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__19734),
            .in2(N__19722),
            .in3(N__19704),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_5_s_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__19701),
            .in2(N__19689),
            .in3(N__19674),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_6_s_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__19671),
            .in2(N__19659),
            .in3(N__19644),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_7_s_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__19641),
            .in2(N__19629),
            .in3(N__19614),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_8_s_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__20055),
            .in2(N__20043),
            .in3(N__20025),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_9_s_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__20022),
            .in2(N__20010),
            .in3(N__19992),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_10_s_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__19989),
            .in2(N__19906),
            .in3(N__19977),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_11_s_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__19897),
            .in2(N__19974),
            .in3(N__19959),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_12_s_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__19956),
            .in2(N__19907),
            .in3(N__19944),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_13_s_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__19901),
            .in2(N__19941),
            .in3(N__19926),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_14_s_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__19923),
            .in2(N__19908),
            .in3(N__19911),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_cry_15_s_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__19905),
            .in2(N__19854),
            .in3(N__19842),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_acc_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_acc_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_16_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164L_LC_1_16_0  (
            .in0(N__20613),
            .in1(N__19839),
            .in2(_gnd_net_),
            .in3(N__20151),
            .lcout(\pwm_generator_inst.un2_threshold_acc_add_1_axb_16_RNI164LZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_17_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_17_2 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_c_RNIFD1K1_LC_1_17_2  (
            .in0(N__21669),
            .in1(N__21686),
            .in2(N__20607),
            .in3(N__21293),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_17_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_RNIRVUI1_LC_1_17_6  (
            .in0(N__22362),
            .in1(N__21351),
            .in2(N__22392),
            .in3(N__21292),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_7_LC_1_18_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_1_18_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_7_LC_1_18_7 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_7_LC_1_18_7  (
            .in0(N__22018),
            .in1(N__20790),
            .in2(N__21939),
            .in3(N__21758),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49211),
            .ce(),
            .sr(N__48542));
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_1_29_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_1_29_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.un7_start_stop_0_a2_LC_1_29_3  (
            .in0(N__48589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23621),
            .lcout(un7_start_stop_0_a2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.N_38_i_i_LC_1_30_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.N_38_i_i_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.N_38_i_i_LC_1_30_0 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \phase_controller_inst1.N_38_i_i_LC_1_30_0  (
            .in0(N__48590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23625),
            .lcout(N_38_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_3  (
            .in0(N__20135),
            .in1(N__20120),
            .in2(_gnd_net_),
            .in3(N__20106),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_2 .LUT_INIT=16'b0011001100000010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_6_2  (
            .in0(N__20408),
            .in1(N__22703),
            .in2(N__22200),
            .in3(N__20286),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_5  (
            .in0(N__20370),
            .in1(N__20355),
            .in2(N__20078),
            .in3(N__20333),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(N__20071),
            .in2(_gnd_net_),
            .in3(N__20254),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_7  (
            .in0(N__20369),
            .in1(N__20354),
            .in2(N__20340),
            .in3(N__20332),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_2  (
            .in0(N__22589),
            .in1(N__22919),
            .in2(N__20988),
            .in3(N__22853),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(\current_shift_inst.PI_CTRL.N_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_7_3 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_7_3  (
            .in0(N__23067),
            .in1(N__20157),
            .in2(N__20310),
            .in3(N__20952),
            .lcout(\current_shift_inst.PI_CTRL.N_153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_7_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_7_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_7_4  (
            .in0(N__20200),
            .in1(N__20219),
            .in2(N__20265),
            .in3(N__20235),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_7_6 .LUT_INIT=16'b1011101110101011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_2_7_6  (
            .in0(N__20229),
            .in1(N__20220),
            .in2(N__20205),
            .in3(N__20184),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_7  (
            .in0(N__23068),
            .in1(_gnd_net_),
            .in2(N__20429),
            .in3(N__22184),
            .lcout(\current_shift_inst.PI_CTRL.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__22656),
            .in2(_gnd_net_),
            .in3(N__22702),
            .lcout(\current_shift_inst.PI_CTRL.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_8_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__22846),
            .in2(_gnd_net_),
            .in3(N__22625),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_8_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_8_6  (
            .in0(N__22918),
            .in1(N__22585),
            .in2(N__20433),
            .in3(N__22887),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(\current_shift_inst.PI_CTRL.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_8_7 .LUT_INIT=16'b0000000011110101;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_8_7  (
            .in0(N__22657),
            .in1(_gnd_net_),
            .in2(N__20412),
            .in3(N__23066),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_2_LC_2_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_2_10_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_2_LC_2_10_1 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_2_LC_2_10_1  (
            .in0(N__21986),
            .in1(N__21852),
            .in2(N__20649),
            .in3(N__21724),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49245),
            .ce(),
            .sr(N__48498));
    defparam \pwm_generator_inst.threshold_ACC_3_LC_2_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_2_10_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_3_LC_2_10_2 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_3_LC_2_10_2  (
            .in0(N__21725),
            .in1(N__21987),
            .in2(N__21911),
            .in3(N__20859),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49245),
            .ce(),
            .sr(N__48498));
    defparam \pwm_generator_inst.threshold_ACC_1_LC_2_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_2_10_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_1_LC_2_10_7 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_1_LC_2_10_7  (
            .in0(N__21985),
            .in1(N__21851),
            .in2(N__20670),
            .in3(N__21723),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49245),
            .ce(),
            .sr(N__48498));
    defparam \pwm_generator_inst.threshold_7_LC_2_11_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_7_LC_2_11_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_7_LC_2_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_7_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20394),
            .lcout(\pwm_generator_inst.thresholdZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49241),
            .ce(),
            .sr(N__48506));
    defparam \pwm_generator_inst.threshold_6_LC_2_12_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_6_LC_2_12_0 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_6_LC_2_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_6_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20382),
            .lcout(\pwm_generator_inst.thresholdZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49237),
            .ce(),
            .sr(N__48516));
    defparam \pwm_generator_inst.threshold_ACC_6_LC_2_12_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_2_12_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_6_LC_2_12_7 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_6_LC_2_12_7  (
            .in0(N__21988),
            .in1(N__21943),
            .in2(N__20814),
            .in3(N__21740),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49237),
            .ce(),
            .sr(N__48516));
    defparam \pwm_generator_inst.threshold_4_LC_2_13_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_4_LC_2_13_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_4_LC_2_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_4_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20376),
            .lcout(\pwm_generator_inst.thresholdZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49233),
            .ce(),
            .sr(N__48522));
    defparam \pwm_generator_inst.threshold_ACC_4_LC_2_13_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_4_LC_2_13_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_4_LC_2_13_6  (
            .in0(N__21741),
            .in1(N__21989),
            .in2(N__21950),
            .in3(N__20841),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49233),
            .ce(),
            .sr(N__48522));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__21251),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TF_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__20529),
            .in2(_gnd_net_),
            .in3(N__20514),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_0_c_RNIE7TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UF_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__20511),
            .in2(_gnd_net_),
            .in3(N__20496),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_1_c_RNIF9UFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVF_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__20493),
            .in2(_gnd_net_),
            .in3(N__20481),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_2_c_RNIGBVFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDO_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__20478),
            .in2(_gnd_net_),
            .in3(N__20472),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_3_c_RNI5LDOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOF_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__38198),
            .in2(N__20469),
            .in3(N__20460),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_4_c_RNI2QOFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQF_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__38200),
            .in2(N__20457),
            .in3(N__20448),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_5_c_RNI4UQFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TF_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__38199),
            .in2(N__20445),
            .in3(N__20436),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_6_c_RNI62TFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_1_9_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__20586),
            .in2(_gnd_net_),
            .in3(N__20580),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_1Z0Z_9 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_9_c_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__20577),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_10_c_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__20571),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_11_c_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__20565),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_12_c_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__20559),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_13_c_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__20553),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_14_c_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__20547),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_15_c_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__20541),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_16_c_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__20535),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_17_c_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__20634),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_18_c_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__20628),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_c_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__20622),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_acc_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_acc_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_acc_cry_19_THRU_LUT4_0_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20616),
            .lcout(\pwm_generator_inst.un3_threshold_acc_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_16_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_c_inv_LC_2_16_5  (
            .in0(N__21527),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20759),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_inv_LC_2_16_6  (
            .in0(N__21687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20600),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_inv_LC_2_16_7  (
            .in0(N__21653),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20690),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_17_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_17_0 .LUT_INIT=16'b1101100001110010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_c_RNIJL5K1_LC_2_17_0  (
            .in0(N__21294),
            .in1(N__21600),
            .in2(N__21207),
            .in3(N__21624),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_inv_LC_2_17_1  (
            .in0(N__20735),
            .in1(N__21591),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_15 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_17_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_17_2 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_RNI91LS1_LC_2_17_2  (
            .in0(N__21296),
            .in1(N__21579),
            .in2(N__20739),
            .in3(N__20736),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_inv_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__21570),
            .in2(_gnd_net_),
            .in3(N__20723),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_16 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_17_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_17_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_c_RNI781K1_LC_2_17_4  (
            .in0(N__20724),
            .in1(N__21558),
            .in2(N__20712),
            .in3(N__21322),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_17_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_inv_LC_2_17_5  (
            .in0(N__21549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20708),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_17 ),
            .ltout(\pwm_generator_inst.un15_threshold_acc_1_axb_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_17_6 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_c_RNIAE4K1_LC_2_17_6  (
            .in0(N__20709),
            .in1(N__21323),
            .in2(N__20697),
            .in3(N__21537),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_17_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_17_7 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_c_RNIHH3K1_LC_2_17_7  (
            .in0(N__21654),
            .in1(N__21633),
            .in2(N__20694),
            .in3(N__21295),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_0_LC_2_18_0  (
            .in0(_gnd_net_),
            .in1(N__20676),
            .in2(N__21335),
            .in3(N__21331),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_18_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_1_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(N__21231),
            .in2(_gnd_net_),
            .in3(N__20658),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_18_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_2_LC_2_18_2  (
            .in0(_gnd_net_),
            .in1(N__20655),
            .in2(_gnd_net_),
            .in3(N__20637),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_18_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_3_LC_2_18_3  (
            .in0(_gnd_net_),
            .in1(N__20865),
            .in2(_gnd_net_),
            .in3(N__20850),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_18_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_4_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(N__20847),
            .in2(_gnd_net_),
            .in3(N__20832),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_18_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_5_LC_2_18_5  (
            .in0(_gnd_net_),
            .in1(N__20829),
            .in2(_gnd_net_),
            .in3(N__20823),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_18_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_18_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_6_LC_2_18_6  (
            .in0(_gnd_net_),
            .in1(N__20820),
            .in2(_gnd_net_),
            .in3(N__20799),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_18_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_18_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_7_LC_2_18_7  (
            .in0(_gnd_net_),
            .in1(N__20796),
            .in2(_gnd_net_),
            .in3(N__20784),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_acc_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_19_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_8_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__20745),
            .in2(_gnd_net_),
            .in3(N__20781),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_2_19_0_),
            .carryout(\pwm_generator_inst.un19_threshold_acc_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_19_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_19_1 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \pwm_generator_inst.threshold_ACC_RNO_0_9_LC_2_19_1  (
            .in0(N__20778),
            .in1(N__21492),
            .in2(N__21336),
            .in3(N__20769),
            .lcout(\pwm_generator_inst.threshold_ACC_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_19_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_19_3 .LUT_INIT=16'b1011100001110100;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_c_RNIDK7K1_LC_2_19_3  (
            .in0(N__21528),
            .in1(N__21327),
            .in2(N__20766),
            .in3(N__21507),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_7_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_7_3  (
            .in0(_gnd_net_),
            .in1(N__22885),
            .in2(_gnd_net_),
            .in3(N__22624),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_3_9_3  (
            .in0(N__22125),
            .in1(N__22212),
            .in2(N__22326),
            .in3(N__22110),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_1_LC_3_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_1_LC_3_10_1 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_1_LC_3_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_1_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20925),
            .lcout(\pwm_generator_inst.thresholdZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49242),
            .ce(),
            .sr(N__48484));
    defparam \pwm_generator_inst.threshold_3_LC_3_10_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_3_LC_3_10_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_3_LC_3_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_3_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20919),
            .lcout(\pwm_generator_inst.thresholdZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49242),
            .ce(),
            .sr(N__48484));
    defparam \pwm_generator_inst.threshold_2_LC_3_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_2_LC_3_10_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_2_LC_3_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_2_LC_3_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20913),
            .lcout(\pwm_generator_inst.thresholdZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49242),
            .ce(),
            .sr(N__48484));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_11_0  (
            .in0(_gnd_net_),
            .in1(N__22077),
            .in2(N__20907),
            .in3(N__22298),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_3_11_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_11_1  (
            .in0(_gnd_net_),
            .in1(N__20898),
            .in2(N__20892),
            .in3(N__22276),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__20883),
            .in2(N__20874),
            .in3(N__22256),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_11_3  (
            .in0(_gnd_net_),
            .in1(N__21102),
            .in2(N__21096),
            .in3(N__22234),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(N__21087),
            .in2(N__21078),
            .in3(N__22555),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_11_5  (
            .in0(_gnd_net_),
            .in1(N__22092),
            .in2(N__21069),
            .in3(N__22534),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_11_6  (
            .in0(_gnd_net_),
            .in1(N__21051),
            .in2(N__21060),
            .in3(N__22513),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_11_7  (
            .in0(N__22492),
            .in1(N__21045),
            .in2(N__21036),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__22029),
            .in2(N__21027),
            .in3(N__22472),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_3_12_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_12_1  (
            .in0(_gnd_net_),
            .in1(N__21018),
            .in2(N__22053),
            .in3(N__22408),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_3_12_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_3_12_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_3_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_3_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21012),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49234),
            .ce(),
            .sr(N__48507));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_3_13_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_3_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_3_13_0  (
            .in0(_gnd_net_),
            .in1(N__22255),
            .in2(_gnd_net_),
            .in3(N__22297),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_3_13_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_3_13_1 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_3_13_1  (
            .in0(N__22556),
            .in1(N__22235),
            .in2(N__21219),
            .in3(N__22277),
            .lcout(\pwm_generator_inst.un1_counterlt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_3_13_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_3_13_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_3_13_4  (
            .in0(N__22493),
            .in1(N__22471),
            .in2(_gnd_net_),
            .in3(N__22409),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto9_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_3_13_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_3_13_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_3_13_5  (
            .in0(N__22515),
            .in1(N__22536),
            .in2(N__21216),
            .in3(N__21213),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_14_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_14_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_c_inv_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(N__21197),
            .in2(_gnd_net_),
            .in3(N__21619),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_0_c_inv_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__21168),
            .in2(_gnd_net_),
            .in3(N__21186),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_0 ),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_1_c_inv_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__21147),
            .in2(_gnd_net_),
            .in3(N__21162),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_2_c_inv_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__21129),
            .in2(_gnd_net_),
            .in3(N__21141),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_3_c_inv_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__21108),
            .in2(_gnd_net_),
            .in3(N__21123),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_4_c_inv_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__21468),
            .in2(_gnd_net_),
            .in3(N__21483),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_5_c_inv_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__21450),
            .in2(_gnd_net_),
            .in3(N__21462),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_6_c_inv_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__21426),
            .in2(_gnd_net_),
            .in3(N__21444),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_7_c_inv_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__21402),
            .in2(_gnd_net_),
            .in3(N__21420),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_8_c_inv_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__21378),
            .in2(_gnd_net_),
            .in3(N__21396),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_8 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_c_inv_LC_3_16_1  (
            .in0(_gnd_net_),
            .in1(N__21357),
            .in2(_gnd_net_),
            .in3(N__21372),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_LUT4_0_LC_3_16_2  (
            .in0(_gnd_net_),
            .in1(N__22357),
            .in2(_gnd_net_),
            .in3(N__21339),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_16_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_RNI3UJI1_LC_3_16_3  (
            .in0(N__21312),
            .in1(N__21255),
            .in2(_gnd_net_),
            .in3(N__21222),
            .lcout(\pwm_generator_inst.un19_threshold_acc_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_16_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_LUT4_0_LC_3_16_4  (
            .in0(_gnd_net_),
            .in1(N__21685),
            .in2(_gnd_net_),
            .in3(N__21657),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_16_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_LUT4_0_LC_3_16_5  (
            .in0(_gnd_net_),
            .in1(N__21649),
            .in2(_gnd_net_),
            .in3(N__21627),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_16_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_LUT4_0_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(N__21620),
            .in2(_gnd_net_),
            .in3(N__21594),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_16_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_LUT4_0_LC_3_16_7  (
            .in0(_gnd_net_),
            .in1(N__21590),
            .in2(_gnd_net_),
            .in3(N__21573),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_LUT4_0_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__21569),
            .in2(_gnd_net_),
            .in3(N__21552),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_LUT4_0_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__21548),
            .in2(_gnd_net_),
            .in3(N__21531),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_LUT4_0_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__21526),
            .in2(_gnd_net_),
            .in3(N__21498),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_acc_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_acc_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_17_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_LUT4_0_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21495),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_18_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_18_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_0_LC_3_18_1 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_0_LC_3_18_1  (
            .in0(N__22008),
            .in1(N__22098),
            .in2(N__21948),
            .in3(N__21761),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49200),
            .ce(),
            .sr(N__48538));
    defparam \pwm_generator_inst.threshold_5_LC_3_18_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_5_LC_3_18_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_5_LC_3_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_5_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22059),
            .lcout(\pwm_generator_inst.thresholdZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49200),
            .ce(),
            .sr(N__48538));
    defparam \pwm_generator_inst.threshold_0_LC_3_18_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_0_LC_3_18_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_0_LC_3_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_0_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22083),
            .lcout(\pwm_generator_inst.thresholdZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49200),
            .ce(),
            .sr(N__48538));
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_18_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_18_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_5_LC_3_18_7 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_5_LC_3_18_7  (
            .in0(N__22009),
            .in1(N__22065),
            .in2(N__21949),
            .in3(N__21762),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49200),
            .ce(),
            .sr(N__48538));
    defparam \pwm_generator_inst.threshold_9_LC_3_19_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_9_LC_3_19_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_9_LC_3_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_9_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22035),
            .lcout(\pwm_generator_inst.thresholdZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49196),
            .ce(),
            .sr(N__48540));
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_19_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_19_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.threshold_ACC_9_LC_3_19_2 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \pwm_generator_inst.threshold_ACC_9_LC_3_19_2  (
            .in0(N__21760),
            .in1(N__22041),
            .in2(N__21951),
            .in3(N__22020),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49196),
            .ce(),
            .sr(N__48540));
    defparam \pwm_generator_inst.threshold_8_LC_3_19_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_8_LC_3_19_4 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_8_LC_3_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.threshold_8_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21693),
            .lcout(\pwm_generator_inst.thresholdZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49196),
            .ce(),
            .sr(N__48540));
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_19_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_19_7 .SEQ_MODE=4'b1011;
    defparam \pwm_generator_inst.threshold_ACC_8_LC_3_19_7 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.threshold_ACC_8_LC_3_19_7  (
            .in0(N__22019),
            .in1(N__21947),
            .in2(N__21771),
            .in3(N__21759),
            .lcout(\pwm_generator_inst.threshold_ACCZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49196),
            .ce(),
            .sr(N__48540));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_9_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_9_2  (
            .in0(N__23033),
            .in1(N__23018),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_9_3  (
            .in0(N__23204),
            .in1(N__23184),
            .in2(N__22215),
            .in3(N__22944),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_10_0  (
            .in0(N__22812),
            .in1(N__22104),
            .in2(N__22797),
            .in3(N__23385),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_10_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_10_1  (
            .in0(N__22332),
            .in1(N__22314),
            .in2(N__22206),
            .in3(N__22305),
            .lcout(\current_shift_inst.PI_CTRL.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_4_10_2  (
            .in0(N__22781),
            .in1(N__22973),
            .in2(N__22992),
            .in3(N__22769),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__22793),
            .in2(_gnd_net_),
            .in3(N__22823),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_10_4  (
            .in0(N__23240),
            .in1(N__23126),
            .in2(N__23228),
            .in3(N__22958),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_10_5  (
            .in0(N__23151),
            .in1(N__22811),
            .in2(N__22119),
            .in3(N__22116),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_10_6  (
            .in0(N__22824),
            .in1(N__23127),
            .in2(N__23019),
            .in3(N__23034),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_10_7  (
            .in0(N__22770),
            .in1(N__22782),
            .in2(N__23229),
            .in3(N__23241),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_11_0  (
            .in0(N__23165),
            .in1(N__23414),
            .in2(N__23403),
            .in3(N__23112),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_11_1  (
            .in0(N__22974),
            .in1(N__23183),
            .in2(N__23205),
            .in3(N__22991),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_11_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_4_11_4  (
            .in0(N__23166),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23111),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_5  (
            .in0(N__23150),
            .in1(N__22943),
            .in2(N__22308),
            .in3(N__22959),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_4_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_4_12_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_4_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_4_12_0  (
            .in0(N__22449),
            .in1(N__22299),
            .in2(_gnd_net_),
            .in3(N__22281),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__49228),
            .ce(),
            .sr(N__48499));
    defparam \pwm_generator_inst.counter_1_LC_4_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_4_12_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_4_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_4_12_1  (
            .in0(N__22443),
            .in1(N__22278),
            .in2(_gnd_net_),
            .in3(N__22260),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__49228),
            .ce(),
            .sr(N__48499));
    defparam \pwm_generator_inst.counter_2_LC_4_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_4_12_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_4_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_4_12_2  (
            .in0(N__22450),
            .in1(N__22257),
            .in2(_gnd_net_),
            .in3(N__22239),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__49228),
            .ce(),
            .sr(N__48499));
    defparam \pwm_generator_inst.counter_3_LC_4_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_4_12_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_4_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_4_12_3  (
            .in0(N__22444),
            .in1(N__22236),
            .in2(_gnd_net_),
            .in3(N__22218),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__49228),
            .ce(),
            .sr(N__48499));
    defparam \pwm_generator_inst.counter_4_LC_4_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_4_12_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_4_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_4_12_4  (
            .in0(N__22451),
            .in1(N__22557),
            .in2(_gnd_net_),
            .in3(N__22539),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__49228),
            .ce(),
            .sr(N__48499));
    defparam \pwm_generator_inst.counter_5_LC_4_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_4_12_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_4_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_4_12_5  (
            .in0(N__22445),
            .in1(N__22535),
            .in2(_gnd_net_),
            .in3(N__22518),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__49228),
            .ce(),
            .sr(N__48499));
    defparam \pwm_generator_inst.counter_6_LC_4_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_4_12_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_4_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_4_12_6  (
            .in0(N__22452),
            .in1(N__22514),
            .in2(_gnd_net_),
            .in3(N__22497),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__49228),
            .ce(),
            .sr(N__48499));
    defparam \pwm_generator_inst.counter_7_LC_4_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_4_12_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_4_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_4_12_7  (
            .in0(N__22446),
            .in1(N__22494),
            .in2(_gnd_net_),
            .in3(N__22476),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__49228),
            .ce(),
            .sr(N__48499));
    defparam \pwm_generator_inst.counter_8_LC_4_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_4_13_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_4_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_4_13_0  (
            .in0(N__22448),
            .in1(N__22473),
            .in2(_gnd_net_),
            .in3(N__22455),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__49222),
            .ce(),
            .sr(N__48508));
    defparam \pwm_generator_inst.counter_9_LC_4_13_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_4_13_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_4_13_1  (
            .in0(N__22410),
            .in1(N__22447),
            .in2(_gnd_net_),
            .in3(N__22413),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49222),
            .ce(),
            .sr(N__48508));
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_4_17_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_4_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_acc_1_cry_10_c_inv_LC_4_17_1  (
            .in0(N__22361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22385),
            .lcout(\pwm_generator_inst.un15_threshold_acc_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_4_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_4_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_4_17_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_4_17_5  (
            .in0(N__33234),
            .in1(N__30126),
            .in2(_gnd_net_),
            .in3(N__33035),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49201),
            .ce(N__32889),
            .sr(N__48533));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_5_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_5_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_5_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22341),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49248),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32460),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49246),
            .ce(),
            .sr(N__48436));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_5_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_5_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_5_7_6  (
            .in0(N__23941),
            .in1(N__28999),
            .in2(N__31907),
            .in3(N__29813),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(N__23337),
            .in2(N__26214),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__49238),
            .ce(),
            .sr(N__48465));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(N__22746),
            .in2(N__32112),
            .in3(N__22725),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__49238),
            .ce(),
            .sr(N__48465));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__28938),
            .in2(N__23328),
            .in3(N__22710),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__49238),
            .ce(),
            .sr(N__48465));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__23316),
            .in2(N__26028),
            .in3(N__22674),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__49238),
            .ce(),
            .sr(N__48465));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__26510),
            .in2(N__23307),
            .in3(N__22635),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__49238),
            .ce(),
            .sr(N__48465));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(N__23358),
            .in2(N__23805),
            .in3(N__22596),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__49238),
            .ce(),
            .sr(N__48465));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__23346),
            .in2(N__26760),
            .in3(N__22926),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__49238),
            .ce(),
            .sr(N__48465));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__23430),
            .in2(N__23733),
            .in3(N__22890),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__49238),
            .ce(),
            .sr(N__48465));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__33366),
            .in2(N__26172),
            .in3(N__22857),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__49235),
            .ce(),
            .sr(N__48471));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__23286),
            .in2(N__26301),
            .in3(N__22827),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__49235),
            .ce(),
            .sr(N__48471));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__27027),
            .in2(N__23277),
            .in3(N__22815),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__49235),
            .ce(),
            .sr(N__48471));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__23295),
            .in2(N__37899),
            .in3(N__22800),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__49235),
            .ce(),
            .sr(N__48471));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__24462),
            .in2(N__32175),
            .in3(N__22785),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__49235),
            .ce(),
            .sr(N__48471));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(N__31908),
            .in2(N__23958),
            .in3(N__22773),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__49235),
            .ce(),
            .sr(N__48471));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(N__23823),
            .in2(N__29004),
            .in3(N__22761),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__49235),
            .ce(),
            .sr(N__48471));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__26357),
            .in2(N__23861),
            .in3(N__23022),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__49235),
            .ce(),
            .sr(N__48471));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__23862),
            .in2(N__23946),
            .in3(N__23001),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__49229),
            .ce(),
            .sr(N__48477));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__32328),
            .in2(N__23892),
            .in3(N__22998),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__49229),
            .ce(),
            .sr(N__48477));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__23866),
            .in2(N__32271),
            .in3(N__22995),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__49229),
            .ce(),
            .sr(N__48477));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__26421),
            .in2(N__23893),
            .in3(N__22977),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__49229),
            .ce(),
            .sr(N__48477));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__23870),
            .in2(N__26850),
            .in3(N__22962),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__49229),
            .ce(),
            .sr(N__48477));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__26898),
            .in2(N__23894),
            .in3(N__22947),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__49229),
            .ce(),
            .sr(N__48477));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__23874),
            .in2(N__31848),
            .in3(N__22929),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__49229),
            .ce(),
            .sr(N__48477));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__29814),
            .in2(N__23895),
            .in3(N__23232),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__49229),
            .ce(),
            .sr(N__48477));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(N__23878),
            .in2(N__26567),
            .in3(N__23208),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__49223),
            .ce(),
            .sr(N__48485));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__44741),
            .in2(N__23896),
            .in3(N__23187),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__49223),
            .ce(),
            .sr(N__48485));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__23882),
            .in2(N__40073),
            .in3(N__23169),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__49223),
            .ce(),
            .sr(N__48485));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__31970),
            .in2(N__23897),
            .in3(N__23154),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__49223),
            .ce(),
            .sr(N__48485));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__23886),
            .in2(N__29223),
            .in3(N__23130),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__49223),
            .ce(),
            .sr(N__48485));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__40314),
            .in2(N__23898),
            .in3(N__23115),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__49223),
            .ce(),
            .sr(N__48485));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__23890),
            .in2(N__26691),
            .in3(N__23103),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__49223),
            .ce(),
            .sr(N__48485));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_12_7  (
            .in0(N__23891),
            .in1(_gnd_net_),
            .in2(N__27357),
            .in3(N__23100),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49223),
            .ce(),
            .sr(N__48485));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_5_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_5_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__29651),
            .in2(_gnd_net_),
            .in3(N__44594),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_5_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_5_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_5_13_5  (
            .in0(N__44595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29597),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_14_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_14_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_5_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_5_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23265),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49213),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_5_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_1_LC_5_16_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_1_LC_5_16_5  (
            .in0(_gnd_net_),
            .in1(N__24560),
            .in2(_gnd_net_),
            .in3(N__23503),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_7_2.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_7_2.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_7_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_7_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23253),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49239),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29805),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_8_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_7_8_0  (
            .in0(N__26166),
            .in1(N__23725),
            .in2(N__26755),
            .in3(N__26291),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_8_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_7_8_1  (
            .in0(N__26509),
            .in1(N__26024),
            .in2(N__23244),
            .in3(N__23801),
            .lcout(\current_shift_inst.PI_CTRL.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_8_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(N__40318),
            .in2(_gnd_net_),
            .in3(N__27022),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_7_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_7_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_7_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32358),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49230),
            .ce(),
            .sr(N__48448));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32685),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49230),
            .ce(),
            .sr(N__48448));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_7_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_7_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_7_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36840),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49230),
            .ce(),
            .sr(N__48448));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_9_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_7_9_4  (
            .in0(N__32436),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49230),
            .ce(),
            .sr(N__48448));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_7_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_7_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_7_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32412),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49230),
            .ce(),
            .sr(N__48448));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_7_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32388),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49230),
            .ce(),
            .sr(N__48448));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32612),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49224),
            .ce(),
            .sr(N__48458));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_7_10_2  (
            .in0(N__33351),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49224),
            .ce(),
            .sr(N__48458));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33447),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49224),
            .ce(),
            .sr(N__48458));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_7_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_7_10_4 .LUT_INIT=16'b0000110011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_7_10_4  (
            .in0(N__27515),
            .in1(N__27355),
            .in2(N__27198),
            .in3(N__24747),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49224),
            .ce(),
            .sr(N__48458));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32654),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49224),
            .ce(),
            .sr(N__48458));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_7_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_7_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26416),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26338),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_7_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_7_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__23418),
            .in2(_gnd_net_),
            .in3(N__23399),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_7_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_7_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23921),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_11_7.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_11_7.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_7_11_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_7_11_7 (
            .in0(N__23373),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49219),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26546),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__23558),
            .in2(_gnd_net_),
            .in3(N__23477),
            .lcout(\phase_controller_inst2.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_7_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_7_13_0 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_7_13_0  (
            .in0(N__35407),
            .in1(N__23987),
            .in2(N__34958),
            .in3(N__23364),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49206),
            .ce(),
            .sr(N__48478));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_13_2 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_7_13_2  (
            .in0(N__24029),
            .in1(N__24052),
            .in2(_gnd_net_),
            .in3(N__24507),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49206),
            .ce(),
            .sr(N__48478));
    defparam \phase_controller_inst2.state_1_LC_7_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_7_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_7_14_2 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst2.state_1_LC_7_14_2  (
            .in0(N__23483),
            .in1(N__23466),
            .in2(N__29961),
            .in3(N__23553),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49202),
            .ce(),
            .sr(N__48486));
    defparam \phase_controller_inst2.state_2_LC_7_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_7_14_4 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \phase_controller_inst2.state_2_LC_7_14_4  (
            .in0(N__29960),
            .in1(N__23465),
            .in2(N__24559),
            .in3(N__23504),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49202),
            .ce(),
            .sr(N__48486));
    defparam \phase_controller_inst2.state_3_LC_7_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_7_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_7_14_6 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \phase_controller_inst2.state_3_LC_7_14_6  (
            .in0(N__23988),
            .in1(N__23505),
            .in2(N__24558),
            .in3(N__31683),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49202),
            .ce(),
            .sr(N__48486));
    defparam \phase_controller_inst2.state_0_LC_7_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_7_14_7 .LUT_INIT=16'b1011101000110000;
    LogicCell40 \phase_controller_inst2.state_0_LC_7_14_7  (
            .in0(N__23554),
            .in1(N__34986),
            .in2(N__24003),
            .in3(N__23484),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49202),
            .ce(),
            .sr(N__48486));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_15_0 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_7_15_0  (
            .in0(N__23643),
            .in1(N__30432),
            .in2(_gnd_net_),
            .in3(N__29982),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_7_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_7_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24054),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__34929),
            .in2(_gnd_net_),
            .in3(N__34957),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_7_15_5  (
            .in0(N__29951),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23464),
            .lcout(\phase_controller_inst2.start_timer_hc_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_15_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_7_15_7  (
            .in0(N__24053),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24030),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_393_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_LC_7_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_7_16_0 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_7_16_0  (
            .in0(N__35400),
            .in1(N__23664),
            .in2(N__23649),
            .in3(N__23658),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49189),
            .ce(),
            .sr(N__48509));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_7_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_7_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_7_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23645),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49189),
            .ce(),
            .sr(N__48509));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_17_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__30433),
            .in2(_gnd_net_),
            .in3(N__23644),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_7_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_7_21_6 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_7_21_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_7_21_6  (
            .in0(N__23608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35396),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49153),
            .ce(),
            .sr(N__48537));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_7_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_7_22_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_7_22_6  (
            .in0(_gnd_net_),
            .in1(N__31717),
            .in2(_gnd_net_),
            .in3(N__31649),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_7_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_7_22_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a2_1_LC_7_22_7  (
            .in0(N__23609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35383),
            .lcout(state_ns_i_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_7_25_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_7_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_7_25_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_7_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23562),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49131),
            .ce(),
            .sr(N__48544));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23520),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49243),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_8_5_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_8_5_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_8_5_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_8_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23511),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49243),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_8_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_8_6_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_8_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24496),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24473),
            .ce(),
            .sr(N__48416));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_7_0  (
            .in0(N__32258),
            .in1(N__31836),
            .in2(N__26420),
            .in3(N__27316),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_8_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_8_7_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_8_7_2  (
            .in0(N__23797),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23729),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_4  (
            .in0(N__23942),
            .in1(N__31886),
            .in2(N__29003),
            .in3(N__29806),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_5  (
            .in0(N__29222),
            .in1(N__23676),
            .in2(N__23697),
            .in3(N__31961),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_8_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_8_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_8_7_6  (
            .in0(N__26553),
            .in1(N__31835),
            .in2(N__32266),
            .in3(N__26411),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_8_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_8_7_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_8_7_7  (
            .in0(N__23682),
            .in1(N__23670),
            .in2(N__23694),
            .in3(N__23691),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_8_8_0  (
            .in0(N__40049),
            .in1(N__44732),
            .in2(N__29221),
            .in3(N__26891),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__26690),
            .in2(_gnd_net_),
            .in3(N__32153),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_8_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_8_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_8_8_3  (
            .in0(N__26831),
            .in1(N__26349),
            .in2(N__32322),
            .in3(N__37881),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_8_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_8_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_8_8_4  (
            .in0(N__26554),
            .in1(N__44733),
            .in2(N__40062),
            .in3(N__26892),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_5  (
            .in0(N__23763),
            .in1(N__23757),
            .in2(N__23751),
            .in3(N__23739),
            .lcout(\current_shift_inst.PI_CTRL.N_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_8_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_8_8_6  (
            .in0(N__26350),
            .in1(N__26832),
            .in2(N__37891),
            .in3(N__32312),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_7  (
            .in0(N__27026),
            .in1(N__40319),
            .in2(N__23748),
            .in3(N__23745),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_8_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_8_9_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_8_9_0  (
            .in0(N__23721),
            .in1(N__44575),
            .in2(N__32613),
            .in3(N__29292),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23720),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_8_9_2 .LUT_INIT=16'b0000000111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_8_9_2  (
            .in0(N__27317),
            .in1(N__27502),
            .in2(N__27176),
            .in3(N__24603),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49225),
            .ce(),
            .sr(N__48437));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_3 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_8_9_3  (
            .in0(N__27501),
            .in1(N__27318),
            .in2(N__24951),
            .in3(N__27132),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49225),
            .ce(),
            .sr(N__48437));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_8_10_2 .LUT_INIT=16'b0000110100011101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_8_10_2  (
            .in0(N__27369),
            .in1(N__27169),
            .in2(N__24855),
            .in3(N__27514),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49220),
            .ce(),
            .sr(N__48449));
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_8_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_8_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32539),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_8_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_8_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_8_10_4  (
            .in0(N__32540),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49220),
            .ce(),
            .sr(N__48449));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_8_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_8_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_8_10_5  (
            .in0(N__29459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44515),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_8_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_8_10_6 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_8_10_6  (
            .in0(N__44516),
            .in1(N__23931),
            .in2(N__23901),
            .in3(N__29445),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_8_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_8_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44517),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49220),
            .ce(),
            .sr(N__48449));
    defparam \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_8_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_8_11_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_8_11_0  (
            .in0(N__23787),
            .in1(N__33347),
            .in2(N__44590),
            .in3(N__29322),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23786),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_8_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_8_11_2 .LUT_INIT=16'b0000000110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_8_11_2  (
            .in0(N__27165),
            .in1(N__27314),
            .in2(N__27524),
            .in3(N__24633),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49214),
            .ce(),
            .sr(N__48459));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_8_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_8_11_3 .LUT_INIT=16'b0010111100101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_8_11_3  (
            .in0(N__27311),
            .in1(N__27167),
            .in2(N__24867),
            .in3(N__27512),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49214),
            .ce(),
            .sr(N__48459));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_8_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_8_11_4 .LUT_INIT=16'b0100010011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_8_11_4  (
            .in0(N__27164),
            .in1(N__27313),
            .in2(N__27523),
            .in3(N__25038),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49214),
            .ce(),
            .sr(N__48459));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_8_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_8_11_5 .LUT_INIT=16'b0010111100101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_8_11_5  (
            .in0(N__27312),
            .in1(N__27168),
            .in2(N__25029),
            .in3(N__27513),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49214),
            .ce(),
            .sr(N__48459));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_8_11_6 .LUT_INIT=16'b0010001000110111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_8_11_6  (
            .in0(N__27166),
            .in1(N__24588),
            .in2(N__27525),
            .in3(N__27315),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49214),
            .ce(),
            .sr(N__48459));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26142),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_8_12_0 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_8_12_0  (
            .in0(N__27516),
            .in1(N__27351),
            .in2(N__24777),
            .in3(N__27160),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49207),
            .ce(),
            .sr(N__48466));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_8_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_8_12_1 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_8_12_1  (
            .in0(N__27350),
            .in1(N__27522),
            .in2(N__27191),
            .in3(N__24900),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49207),
            .ce(),
            .sr(N__48466));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_8_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_8_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_8_12_2 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_8_12_2  (
            .in0(N__27518),
            .in1(N__27353),
            .in2(N__24879),
            .in3(N__27162),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49207),
            .ce(),
            .sr(N__48466));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_8_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_8_12_3 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_8_12_3  (
            .in0(N__27349),
            .in1(N__27521),
            .in2(N__27190),
            .in3(N__24924),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49207),
            .ce(),
            .sr(N__48466));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_8_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_8_12_4 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_8_12_4  (
            .in0(N__27517),
            .in1(N__27352),
            .in2(N__24936),
            .in3(N__27161),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49207),
            .ce(),
            .sr(N__48466));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_8_12_5 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_8_12_5  (
            .in0(N__27348),
            .in1(N__27520),
            .in2(N__27189),
            .in3(N__24984),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49207),
            .ce(),
            .sr(N__48466));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_6 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_8_12_6  (
            .in0(N__27519),
            .in1(N__27354),
            .in2(N__25002),
            .in3(N__27163),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49207),
            .ce(),
            .sr(N__48466));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_13_0 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_8_13_0  (
            .in0(N__24503),
            .in1(N__24051),
            .in2(_gnd_net_),
            .in3(N__24028),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_394_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_8_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_8_14_0 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_8_14_0  (
            .in0(N__31128),
            .in1(N__30786),
            .in2(N__29091),
            .in3(N__47699),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_8_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_8_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__34985),
            .in2(_gnd_net_),
            .in3(N__23999),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_8_15_0  (
            .in0(N__24267),
            .in1(N__28042),
            .in2(_gnd_net_),
            .in3(N__23976),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__49190),
            .ce(N__24145),
            .sr(N__48487));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_8_15_1  (
            .in0(N__24241),
            .in1(N__27989),
            .in2(_gnd_net_),
            .in3(N__23973),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__49190),
            .ce(N__24145),
            .sr(N__48487));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_8_15_2  (
            .in0(N__24268),
            .in1(N__27937),
            .in2(_gnd_net_),
            .in3(N__23970),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__49190),
            .ce(N__24145),
            .sr(N__48487));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_8_15_3  (
            .in0(N__24242),
            .in1(N__27878),
            .in2(_gnd_net_),
            .in3(N__23967),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__49190),
            .ce(N__24145),
            .sr(N__48487));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_8_15_4  (
            .in0(N__24269),
            .in1(N__27824),
            .in2(_gnd_net_),
            .in3(N__23964),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__49190),
            .ce(N__24145),
            .sr(N__48487));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_8_15_5  (
            .in0(N__24243),
            .in1(N__28336),
            .in2(_gnd_net_),
            .in3(N__23961),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__49190),
            .ce(N__24145),
            .sr(N__48487));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_8_15_6  (
            .in0(N__24270),
            .in1(N__28310),
            .in2(_gnd_net_),
            .in3(N__24081),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__49190),
            .ce(N__24145),
            .sr(N__48487));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_8_15_7  (
            .in0(N__24244),
            .in1(N__28291),
            .in2(_gnd_net_),
            .in3(N__24078),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__49190),
            .ce(N__24145),
            .sr(N__48487));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_8_16_0  (
            .in0(N__24248),
            .in1(N__28255),
            .in2(_gnd_net_),
            .in3(N__24075),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__49182),
            .ce(N__24144),
            .sr(N__48500));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_8_16_1  (
            .in0(N__24252),
            .in1(N__28225),
            .in2(_gnd_net_),
            .in3(N__24072),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__49182),
            .ce(N__24144),
            .sr(N__48500));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_8_16_2  (
            .in0(N__24245),
            .in1(N__28189),
            .in2(_gnd_net_),
            .in3(N__24069),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__49182),
            .ce(N__24144),
            .sr(N__48500));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_8_16_3  (
            .in0(N__24249),
            .in1(N__28154),
            .in2(_gnd_net_),
            .in3(N__24066),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__49182),
            .ce(N__24144),
            .sr(N__48500));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_8_16_4  (
            .in0(N__24246),
            .in1(N__28130),
            .in2(_gnd_net_),
            .in3(N__24063),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__49182),
            .ce(N__24144),
            .sr(N__48500));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_16_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_8_16_5  (
            .in0(N__24250),
            .in1(N__28100),
            .in2(_gnd_net_),
            .in3(N__24060),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__49182),
            .ce(N__24144),
            .sr(N__48500));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_16_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_16_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_8_16_6  (
            .in0(N__24247),
            .in1(N__28571),
            .in2(_gnd_net_),
            .in3(N__24057),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__49182),
            .ce(N__24144),
            .sr(N__48500));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_16_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_8_16_7  (
            .in0(N__24251),
            .in1(N__28537),
            .in2(_gnd_net_),
            .in3(N__24108),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__49182),
            .ce(N__24144),
            .sr(N__48500));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_8_17_0  (
            .in0(N__24263),
            .in1(N__28507),
            .in2(_gnd_net_),
            .in3(N__24105),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__49174),
            .ce(N__24146),
            .sr(N__48510));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_8_17_1  (
            .in0(N__24253),
            .in1(N__28480),
            .in2(_gnd_net_),
            .in3(N__24102),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__49174),
            .ce(N__24146),
            .sr(N__48510));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_8_17_2  (
            .in0(N__24264),
            .in1(N__28459),
            .in2(_gnd_net_),
            .in3(N__24099),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__49174),
            .ce(N__24146),
            .sr(N__48510));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_8_17_3  (
            .in0(N__24254),
            .in1(N__28429),
            .in2(_gnd_net_),
            .in3(N__24096),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__49174),
            .ce(N__24146),
            .sr(N__48510));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_8_17_4  (
            .in0(N__24265),
            .in1(N__28394),
            .in2(_gnd_net_),
            .in3(N__24093),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__49174),
            .ce(N__24146),
            .sr(N__48510));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_8_17_5  (
            .in0(N__24255),
            .in1(N__28366),
            .in2(_gnd_net_),
            .in3(N__24090),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__49174),
            .ce(N__24146),
            .sr(N__48510));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_8_17_6  (
            .in0(N__24266),
            .in1(N__28883),
            .in2(_gnd_net_),
            .in3(N__24087),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__49174),
            .ce(N__24146),
            .sr(N__48510));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_8_17_7  (
            .in0(N__24256),
            .in1(N__28859),
            .in2(_gnd_net_),
            .in3(N__24084),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__49174),
            .ce(N__24146),
            .sr(N__48510));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_8_18_0  (
            .in0(N__24257),
            .in1(N__28828),
            .in2(_gnd_net_),
            .in3(N__24285),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__49167),
            .ce(N__24150),
            .sr(N__48517));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_8_18_1  (
            .in0(N__24261),
            .in1(N__28775),
            .in2(_gnd_net_),
            .in3(N__24282),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__49167),
            .ce(N__24150),
            .sr(N__48517));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_8_18_2  (
            .in0(N__24258),
            .in1(N__28735),
            .in2(_gnd_net_),
            .in3(N__24279),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__49167),
            .ce(N__24150),
            .sr(N__48517));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_8_18_3  (
            .in0(N__24262),
            .in1(N__28658),
            .in2(_gnd_net_),
            .in3(N__24276),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__49167),
            .ce(N__24150),
            .sr(N__48517));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_8_18_4  (
            .in0(N__24259),
            .in1(N__28709),
            .in2(_gnd_net_),
            .in3(N__24273),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__49167),
            .ce(N__24150),
            .sr(N__48517));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_18_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_8_18_5  (
            .in0(N__28688),
            .in1(N__24260),
            .in2(_gnd_net_),
            .in3(N__24153),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49167),
            .ce(N__24150),
            .sr(N__48517));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28053),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49159),
            .ce(N__28620),
            .sr(N__48523));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3 .LUT_INIT=16'b1101000011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_8_20_3  (
            .in0(N__25689),
            .in1(N__31558),
            .in2(N__31722),
            .in3(N__24339),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49154),
            .ce(),
            .sr(N__48528));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_21_4 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_8_21_4  (
            .in0(N__24334),
            .in1(N__24351),
            .in2(N__25203),
            .in3(N__32765),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49148),
            .ce(),
            .sr(N__48534));
    defparam \phase_controller_inst1.stoper_hc.running_LC_8_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_8_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_8_21_7 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_8_21_7  (
            .in0(N__31718),
            .in1(N__25688),
            .in2(N__24366),
            .in3(N__24335),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49148),
            .ce(),
            .sr(N__48534));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_8_22_0  (
            .in0(_gnd_net_),
            .in1(N__24332),
            .in2(_gnd_net_),
            .in3(N__24350),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_22_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_8_22_1  (
            .in0(N__31706),
            .in1(N__24362),
            .in2(_gnd_net_),
            .in3(N__31648),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_8_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_8_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_8_22_2 .LUT_INIT=16'b1111111100111011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_8_22_2  (
            .in0(N__25704),
            .in1(N__31707),
            .in2(N__25635),
            .in3(N__25664),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_8_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_8_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_8_22_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_8_22_3  (
            .in0(N__24333),
            .in1(_gnd_net_),
            .in2(N__24312),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_23_0  (
            .in0(_gnd_net_),
            .in1(N__25202),
            .in2(N__24309),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_23_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_23_1  (
            .in0(N__32758),
            .in1(N__25155),
            .in2(_gnd_net_),
            .in3(N__24300),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49137),
            .ce(),
            .sr(N__48539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_23_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_23_2  (
            .in0(N__32762),
            .in1(N__24297),
            .in2(N__25425),
            .in3(N__24291),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49137),
            .ce(),
            .sr(N__48539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_23_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_23_3  (
            .in0(N__32759),
            .in1(N__25389),
            .in2(_gnd_net_),
            .in3(N__24288),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49137),
            .ce(),
            .sr(N__48539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_23_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_23_4  (
            .in0(N__32763),
            .in1(N__25368),
            .in2(_gnd_net_),
            .in3(N__24393),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49137),
            .ce(),
            .sr(N__48539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_23_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_23_5  (
            .in0(N__32760),
            .in1(N__25320),
            .in2(_gnd_net_),
            .in3(N__24390),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49137),
            .ce(),
            .sr(N__48539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_23_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_23_6  (
            .in0(N__32764),
            .in1(N__25284),
            .in2(_gnd_net_),
            .in3(N__24387),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49137),
            .ce(),
            .sr(N__48539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_23_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_23_7  (
            .in0(N__32761),
            .in1(N__25263),
            .in2(_gnd_net_),
            .in3(N__24384),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49137),
            .ce(),
            .sr(N__48539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_24_0  (
            .in0(N__32866),
            .in1(N__25233),
            .in2(_gnd_net_),
            .in3(N__24381),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_24_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49132),
            .ce(),
            .sr(N__48541));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_24_1  (
            .in0(N__32851),
            .in1(N__25605),
            .in2(_gnd_net_),
            .in3(N__24378),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49132),
            .ce(),
            .sr(N__48541));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_24_2  (
            .in0(N__32863),
            .in1(N__25572),
            .in2(_gnd_net_),
            .in3(N__24375),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49132),
            .ce(),
            .sr(N__48541));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_24_3  (
            .in0(N__32852),
            .in1(N__25542),
            .in2(_gnd_net_),
            .in3(N__24372),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49132),
            .ce(),
            .sr(N__48541));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_24_4  (
            .in0(N__32864),
            .in1(N__25515),
            .in2(_gnd_net_),
            .in3(N__24369),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49132),
            .ce(),
            .sr(N__48541));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_24_5  (
            .in0(N__32853),
            .in1(N__25485),
            .in2(_gnd_net_),
            .in3(N__24420),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49132),
            .ce(),
            .sr(N__48541));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_24_6  (
            .in0(N__32865),
            .in1(N__25452),
            .in2(_gnd_net_),
            .in3(N__24417),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49132),
            .ce(),
            .sr(N__48541));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_24_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_24_7  (
            .in0(N__32854),
            .in1(N__25791),
            .in2(_gnd_net_),
            .in3(N__24414),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49132),
            .ce(),
            .sr(N__48541));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_25_0  (
            .in0(N__32855),
            .in1(N__25824),
            .in2(_gnd_net_),
            .in3(N__24411),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_8_25_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49125),
            .ce(),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_25_1  (
            .in0(N__32859),
            .in1(N__25896),
            .in2(_gnd_net_),
            .in3(N__24408),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49125),
            .ce(),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_25_2  (
            .in0(N__32856),
            .in1(N__25880),
            .in2(_gnd_net_),
            .in3(N__24405),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49125),
            .ce(),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_25_3  (
            .in0(N__32860),
            .in1(N__25842),
            .in2(_gnd_net_),
            .in3(N__24402),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49125),
            .ce(),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_25_4  (
            .in0(N__32857),
            .in1(N__25854),
            .in2(_gnd_net_),
            .in3(N__24399),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49125),
            .ce(),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_25_5  (
            .in0(N__32861),
            .in1(N__25755),
            .in2(_gnd_net_),
            .in3(N__24396),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49125),
            .ce(),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_25_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_25_6  (
            .in0(N__32858),
            .in1(N__25767),
            .in2(_gnd_net_),
            .in3(N__24447),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49125),
            .ce(),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_25_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_25_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_25_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_25_7  (
            .in0(N__32862),
            .in1(N__25929),
            .in2(_gnd_net_),
            .in3(N__24444),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49125),
            .ce(),
            .sr(N__48543));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_26_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_26_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_26_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_26_0  (
            .in0(N__32844),
            .in1(N__25941),
            .in2(_gnd_net_),
            .in3(N__24441),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_8_26_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49121),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_26_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_26_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_26_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_26_1  (
            .in0(N__32848),
            .in1(N__25737),
            .in2(_gnd_net_),
            .in3(N__24438),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49121),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_26_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_26_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_26_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_26_2  (
            .in0(N__32845),
            .in1(N__25725),
            .in2(_gnd_net_),
            .in3(N__24435),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49121),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_26_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_26_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_26_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_26_3  (
            .in0(N__32849),
            .in1(N__26094),
            .in2(_gnd_net_),
            .in3(N__24432),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49121),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_26_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_26_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_26_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_26_4  (
            .in0(N__32846),
            .in1(N__26106),
            .in2(_gnd_net_),
            .in3(N__24429),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49121),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_26_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_26_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_26_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_26_5  (
            .in0(N__32850),
            .in1(N__25631),
            .in2(_gnd_net_),
            .in3(N__24426),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49121),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_26_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_26_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_26_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_26_6  (
            .in0(N__32847),
            .in1(N__25663),
            .in2(_gnd_net_),
            .in3(N__24423),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49121),
            .ce(),
            .sr(N__48545));
    defparam \phase_controller_inst2.S1_LC_8_30_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_8_30_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_8_30_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_8_30_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24567),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49112),
            .ce(),
            .sr(N__48546));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_5_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26499),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_5_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_5_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_5_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_9_5_1 (
            .in0(N__24516),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49240),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_9_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_9_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_9_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24495),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24474),
            .ce(),
            .sr(N__48408));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_9_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_9_7_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_9_7_0 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_9_7_0  (
            .in0(N__27370),
            .in1(N__27477),
            .in2(N__27177),
            .in3(N__24669),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49231),
            .ce(),
            .sr(N__48417));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_9_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_9_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32573),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49231),
            .ce(),
            .sr(N__48417));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_9_7_3 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_9_7_3  (
            .in0(N__27473),
            .in1(N__27137),
            .in2(_gnd_net_),
            .in3(N__24579),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49231),
            .ce(),
            .sr(N__48417));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_7_4 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_9_7_4  (
            .in0(N__27133),
            .in1(N__27476),
            .in2(_gnd_net_),
            .in3(N__24714),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49231),
            .ce(),
            .sr(N__48417));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_9_7_5 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_9_7_5  (
            .in0(N__27474),
            .in1(N__27371),
            .in2(N__24732),
            .in3(N__27138),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49231),
            .ce(),
            .sr(N__48417));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_9_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_9_7_7 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_9_7_7  (
            .in0(N__27475),
            .in1(N__27372),
            .in2(N__24966),
            .in3(N__27139),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49231),
            .ce(),
            .sr(N__48417));
    defparam \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_9_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_9_8_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_9_8_0  (
            .in0(N__26013),
            .in1(N__32655),
            .in2(N__44598),
            .in3(N__29103),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26012),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_2 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_9_8_2  (
            .in0(N__27126),
            .in1(N__27438),
            .in2(_gnd_net_),
            .in3(N__24687),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49226),
            .ce(),
            .sr(N__48422));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_9_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_9_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_9_8_3 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_9_8_3  (
            .in0(N__27434),
            .in1(N__27360),
            .in2(N__24840),
            .in3(N__27127),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49226),
            .ce(),
            .sr(N__48422));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_8_4 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_9_8_4  (
            .in0(N__27358),
            .in1(N__27436),
            .in2(N__27174),
            .in3(N__24825),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49226),
            .ce(),
            .sr(N__48422));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_8_5 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_9_8_5  (
            .in0(N__27435),
            .in1(N__27361),
            .in2(N__24813),
            .in3(N__27128),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49226),
            .ce(),
            .sr(N__48422));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_9_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_9_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_9_8_6 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_9_8_6  (
            .in0(N__27359),
            .in1(N__27437),
            .in2(N__27175),
            .in3(N__24798),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49226),
            .ce(),
            .sr(N__48422));
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__26636),
            .in2(N__26640),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_9_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__26244),
            .in2(N__26235),
            .in3(N__24570),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_9_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__26220),
            .in2(N__32067),
            .in3(N__24717),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_9_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_9_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__28902),
            .in2(N__26442),
            .in3(N__24705),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_9_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_9_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__24702),
            .in2(N__24696),
            .in3(N__24681),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__24678),
            .in2(N__26466),
            .in3(N__24660),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__24657),
            .in2(N__24645),
            .in3(N__24624),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__26781),
            .in2(N__26796),
            .in3(N__24621),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__24618),
            .in2(N__24612),
            .in3(N__24597),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__24594),
            .in2(N__26121),
            .in3(N__24582),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__26073),
            .in2(N__26253),
            .in3(N__24846),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__26112),
            .in2(N__26181),
            .in3(N__24843),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__37848),
            .in2(N__26430),
            .in3(N__24828),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__32124),
            .in2(N__26625),
            .in3(N__24816),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__31860),
            .in2(N__26313),
            .in3(N__24801),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__28950),
            .in2(N__26649),
            .in3(N__24789),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__24786),
            .in2(N__26322),
            .in3(N__24768),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__24765),
            .in2(N__24756),
            .in3(N__24735),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__32283),
            .in2(N__26616),
            .in3(N__24987),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__32220),
            .in2(N__26586),
            .in3(N__24978),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__24975),
            .in2(N__26373),
            .in3(N__24954),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__25959),
            .in2(N__26805),
            .in3(N__24939),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__26859),
            .in2(N__26595),
            .in3(N__24927),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__31800),
            .in2(N__26607),
            .in3(N__24918),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__24915),
            .in2(N__29754),
            .in3(N__24891),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__24888),
            .in2(N__26520),
            .in3(N__24870),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__44694),
            .in2(N__29838),
            .in3(N__24858),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__40017),
            .in2(N__26577),
            .in3(N__25032),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__31923),
            .in2(N__29547),
            .in3(N__25017),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__29884),
            .in2(N__29169),
            .in3(N__25014),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__29886),
            .in2(N__40278),
            .in3(N__25011),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__29885),
            .in2(N__26457),
            .in3(N__25008),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_9_13_0  (
            .in0(N__27277),
            .in1(N__44565),
            .in2(_gnd_net_),
            .in3(N__25005),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_9_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_9_13_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__24993),
            .in2(_gnd_net_),
            .in3(N__47691),
            .lcout(elapsed_time_ns_1_RNIRB3CP1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_9_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_9_14_0 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_9_14_0  (
            .in0(N__31105),
            .in1(N__28026),
            .in2(N__30255),
            .in3(N__30155),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_9_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_9_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_9_14_2 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_9_14_2  (
            .in0(N__33293),
            .in1(N__30154),
            .in2(N__29676),
            .in3(N__32997),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49191),
            .ce(N__32900),
            .sr(N__48472));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_9_14_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_9_14_3 .LUT_INIT=16'b1111111111100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_9_14_3  (
            .in0(N__30001),
            .in1(N__31106),
            .in2(N__27864),
            .in3(N__47703),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_9_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_9_14_4 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_9_14_4  (
            .in0(N__30251),
            .in1(_gnd_net_),
            .in2(N__25047),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIUE3CP1_0_6),
            .ltout(elapsed_time_ns_1_RNIUE3CP1_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_9_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_9_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_9_14_5 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_9_14_5  (
            .in0(N__32996),
            .in1(N__33229),
            .in2(N__25044),
            .in3(N__33294),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49191),
            .ce(N__32900),
            .sr(N__48472));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_14_7 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_9_14_7  (
            .in0(N__32995),
            .in1(N__27569),
            .in2(N__33309),
            .in3(N__33230),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49191),
            .ce(N__32900),
            .sr(N__48472));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_15_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_9_15_1  (
            .in0(N__33202),
            .in1(N__30057),
            .in2(N__31400),
            .in3(N__27628),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49183),
            .ce(N__32901),
            .sr(N__48479));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_9_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_9_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_9_15_2 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_9_15_2  (
            .in0(N__27585),
            .in1(N__30195),
            .in2(N__27597),
            .in3(N__33314),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49183),
            .ce(N__32901),
            .sr(N__48479));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_9_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_9_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_9_15_3 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_9_15_3  (
            .in0(N__33203),
            .in1(N__28083),
            .in2(N__33315),
            .in3(N__33003),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49183),
            .ce(N__32901),
            .sr(N__48479));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_9_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_9_16_0 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_9_16_0  (
            .in0(N__30762),
            .in1(N__31093),
            .in2(N__25106),
            .in3(N__47702),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_9_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_9_16_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25041),
            .in3(N__30231),
            .lcout(elapsed_time_ns_1_RNIFFC6P1_0_16),
            .ltout(elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_9_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_9_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_9_16_2 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_9_16_2  (
            .in0(N__33240),
            .in1(_gnd_net_),
            .in2(N__25074),
            .in3(N__31371),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49175),
            .ce(N__34507),
            .sr(N__48488));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_16_3 .LUT_INIT=16'b1000111010101111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_9_16_3  (
            .in0(N__25061),
            .in1(N__25070),
            .in2(N__34038),
            .in3(N__34064),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_16_4 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_16_4  (
            .in0(N__25071),
            .in1(N__25062),
            .in2(N__34065),
            .in3(N__34037),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_9_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_9_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_9_16_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_9_16_5  (
            .in0(N__31370),
            .in1(N__33242),
            .in2(_gnd_net_),
            .in3(N__29090),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49175),
            .ce(N__34507),
            .sr(N__48488));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_16_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_9_16_6  (
            .in0(N__33241),
            .in1(N__30945),
            .in2(_gnd_net_),
            .in3(N__31372),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49175),
            .ce(N__34507),
            .sr(N__48488));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_16_7 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_16_7  (
            .in0(N__31272),
            .in1(N__34253),
            .in2(N__34224),
            .in3(N__31247),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_9_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_9_17_0 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_9_17_0  (
            .in0(N__31043),
            .in1(N__30655),
            .in2(N__27565),
            .in3(N__27977),
            .lcout(elapsed_time_ns_1_RNILGKEE1_0_4),
            .ltout(elapsed_time_ns_1_RNILGKEE1_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_9_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_9_17_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_9_17_1  (
            .in0(N__30938),
            .in1(N__28077),
            .in2(N__25053),
            .in3(N__31290),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_9_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_9_17_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_9_17_2  (
            .in0(N__29064),
            .in1(_gnd_net_),
            .in2(N__25050),
            .in3(N__25104),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_9_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_9_17_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_9_17_3  (
            .in0(N__25105),
            .in1(N__29065),
            .in2(N__30949),
            .in3(N__31291),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_17_4 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__27734),
            .in2(N__25134),
            .in3(N__30051),
            .lcout(\phase_controller_inst1.stoper_hc.N_316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_9_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_9_17_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_9_17_5  (
            .in0(N__48588),
            .in1(N__27778),
            .in2(_gnd_net_),
            .in3(N__47633),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_342_i ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_342_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_9_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_9_17_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25131),
            .in3(N__25125),
            .lcout(elapsed_time_ns_1_RNIHHC6P1_0_18),
            .ltout(elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_9_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_9_17_7 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_9_17_7  (
            .in0(N__30743),
            .in1(N__31042),
            .in2(N__25128),
            .in3(N__47634),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_9_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_9_18_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__25119),
            .in2(_gnd_net_),
            .in3(N__30238),
            .lcout(elapsed_time_ns_1_RNIGGC6P1_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_18_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_9_18_5  (
            .in0(N__31429),
            .in1(N__33121),
            .in2(_gnd_net_),
            .in3(N__25107),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49160),
            .ce(N__32896),
            .sr(N__48511));
    defparam \phase_controller_inst1.stoper_hc.N_267_i_1_LC_9_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.N_267_i_1_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.N_267_i_1_LC_9_19_1 .LUT_INIT=16'b0011001100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.N_267_i_1_LC_9_19_1  (
            .in0(N__27754),
            .in1(N__27629),
            .in2(N__30330),
            .in3(N__30064),
            .lcout(\phase_controller_inst1.stoper_hc.N_267_iZ0Z_1 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_267_iZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_9_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_9_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_9_19_2 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_9_19_2  (
            .in0(N__26922),
            .in1(N__33120),
            .in2(N__25077),
            .in3(N__31425),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49155),
            .ce(N__34575),
            .sr(N__48518));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_9_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_9_19_3 .LUT_INIT=16'b1111111111100100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_9_19_3  (
            .in0(N__31124),
            .in1(N__26923),
            .in2(N__29741),
            .in3(N__47698),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_9_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_9_19_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25212),
            .in3(N__30252),
            .lcout(elapsed_time_ns_1_RNI1I3CP1_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_9_19_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_9_19_5  (
            .in0(N__33119),
            .in1(N__30065),
            .in2(N__31441),
            .in3(N__27630),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49155),
            .ce(N__34575),
            .sr(N__48518));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_9_19_7 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_9_19_7  (
            .in0(N__33118),
            .in1(N__27758),
            .in2(N__31440),
            .in3(N__31479),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49155),
            .ce(N__34575),
            .sr(N__48518));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_5 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_9_20_5  (
            .in0(N__33239),
            .in1(N__25209),
            .in2(N__31442),
            .in3(N__26921),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49149),
            .ce(N__32897),
            .sr(N__48524));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_21_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_9_21_1  (
            .in0(N__31437),
            .in1(N__33237),
            .in2(N__30501),
            .in3(N__31494),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49142),
            .ce(N__32898),
            .sr(N__48529));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_21_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_9_21_2  (
            .in0(N__33235),
            .in1(N__31541),
            .in2(N__31504),
            .in3(N__31439),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49142),
            .ce(N__32898),
            .sr(N__48529));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_9_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_9_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_9_21_3 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_9_21_3  (
            .in0(N__31438),
            .in1(N__33238),
            .in2(N__27762),
            .in3(N__31495),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49142),
            .ce(N__32898),
            .sr(N__48529));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_9_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_9_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_9_21_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_9_21_5  (
            .in0(N__30539),
            .in1(N__33236),
            .in2(N__31443),
            .in3(N__31493),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49142),
            .ce(N__32898),
            .sr(N__48529));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_9_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_9_22_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_9_22_0  (
            .in0(N__25201),
            .in1(N__25176),
            .in2(N__25164),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_9_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_9_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(N__32919),
            .in2(N__25143),
            .in3(N__25154),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_9_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_9_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_9_22_2  (
            .in0(_gnd_net_),
            .in1(N__25434),
            .in2(N__25410),
            .in3(N__25421),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_9_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_9_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(N__25401),
            .in2(N__25377),
            .in3(N__25388),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_9_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_9_22_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_9_22_4  (
            .in0(N__25367),
            .in1(N__25356),
            .in2(N__25347),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_9_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_9_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__25335),
            .in2(N__25308),
            .in3(N__25319),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_9_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_9_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__25299),
            .in2(N__25272),
            .in3(N__25283),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_9_22_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_9_22_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_9_22_7  (
            .in0(N__25262),
            .in1(N__29010),
            .in2(N__25251),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_9_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_9_23_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_9_23_0  (
            .in0(_gnd_net_),
            .in1(N__25242),
            .in2(N__25221),
            .in3(N__25232),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_9_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_9_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_9_23_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_9_23_1  (
            .in0(_gnd_net_),
            .in1(N__29031),
            .in2(N__25593),
            .in3(N__25604),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_9_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_9_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_9_23_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_9_23_2  (
            .in0(_gnd_net_),
            .in1(N__25560),
            .in2(N__25584),
            .in3(N__25571),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_9_23_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_9_23_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_9_23_3  (
            .in0(_gnd_net_),
            .in1(N__25530),
            .in2(N__25554),
            .in3(N__25541),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_9_23_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_9_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_9_23_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__25524),
            .in2(N__25503),
            .in3(N__25514),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_9_23_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_9_23_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(N__25494),
            .in2(N__25473),
            .in3(N__25484),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_9_23_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_9_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_9_23_6  (
            .in0(_gnd_net_),
            .in1(N__25440),
            .in2(N__25464),
            .in3(N__25451),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_9_23_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_9_23_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_9_23_7  (
            .in0(_gnd_net_),
            .in1(N__25776),
            .in2(N__25911),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_9_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_9_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__25947),
            .in2(N__25863),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_9_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_9_24_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__25830),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_9_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_9_24_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_9_24_2  (
            .in0(_gnd_net_),
            .in1(N__25743),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_9_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_9_24_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__25917),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_9_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_9_24_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(N__25713),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_9_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_9_24_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(N__26082),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_9_24_6  (
            .in0(_gnd_net_),
            .in1(N__25611),
            .in2(N__25668),
            .in3(N__25695),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25692),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_9_25_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_9_25_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_9_25_0  (
            .in0(_gnd_net_),
            .in1(N__25659),
            .in2(_gnd_net_),
            .in3(N__25630),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_25_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_25_1 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_25_1  (
            .in0(N__25894),
            .in1(N__25876),
            .in2(N__29025),
            .in3(N__28599),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_25_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_25_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__25940),
            .in2(_gnd_net_),
            .in3(N__25928),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_25_3 .LUT_INIT=16'b0111001100010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_25_3  (
            .in0(N__25790),
            .in1(N__25823),
            .in2(N__25809),
            .in3(N__29045),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_25_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_25_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_25_4  (
            .in0(N__28598),
            .in1(N__25895),
            .in2(N__25881),
            .in3(N__29024),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_9_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_9_25_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_9_25_5  (
            .in0(_gnd_net_),
            .in1(N__25853),
            .in2(_gnd_net_),
            .in3(N__25841),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_9_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_9_25_6 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_9_25_6  (
            .in0(N__25822),
            .in1(N__25808),
            .in2(N__29046),
            .in3(N__25789),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_25_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_25_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_25_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_25_7  (
            .in0(_gnd_net_),
            .in1(N__25766),
            .in2(_gnd_net_),
            .in3(N__25754),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_9_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_9_26_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_9_26_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_9_26_2  (
            .in0(_gnd_net_),
            .in1(N__25736),
            .in2(_gnd_net_),
            .in3(N__25724),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_9_26_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_9_26_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_9_26_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_9_26_6  (
            .in0(_gnd_net_),
            .in1(N__26105),
            .in2(_gnd_net_),
            .in3(N__26093),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26299),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_10_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_10_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__29389),
            .in2(_gnd_net_),
            .in3(N__44586),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_10_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_10_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_10_7_2  (
            .in0(N__26683),
            .in1(N__31969),
            .in2(N__32167),
            .in3(N__27356),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_10_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_10_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_10_7_3  (
            .in0(N__26061),
            .in1(N__26052),
            .in2(N__26043),
            .in3(N__25989),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_10_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_10_7_4 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_10_7_4  (
            .in0(N__26167),
            .in1(N__26040),
            .in2(N__26759),
            .in3(N__26300),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_10_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_10_7_5 .LUT_INIT=16'b1111001011110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_10_7_5  (
            .in0(N__26187),
            .in1(N__26492),
            .in2(N__26031),
            .in3(N__26020),
            .lcout(\current_shift_inst.PI_CTRL.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_10_7_6 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_10_7_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_10_7_6  (
            .in0(N__48583),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_10_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_10_7_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_10_7_7  (
            .in0(N__26845),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_10_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_10_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32383),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_10_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_10_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26200),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_0 ),
            .ltout(\current_shift_inst.PI_CTRL.integrator_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_10_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_10_8_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_10_8_3  (
            .in0(N__32384),
            .in1(N__44535),
            .in2(N__26238),
            .in3(N__29124),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_8_4 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_10_8_4  (
            .in0(N__27170),
            .in1(N__27439),
            .in2(_gnd_net_),
            .in3(N__26226),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49215),
            .ce(),
            .sr(N__48412));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32091),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_10_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_10_8_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_10_8_6  (
            .in0(N__32092),
            .in1(N__28929),
            .in2(_gnd_net_),
            .in3(N__26201),
            .lcout(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_10_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_10_9_0 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_10_9_0  (
            .in0(N__32508),
            .in1(N__27009),
            .in2(N__44597),
            .in3(N__29244),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_10_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_10_9_1 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_10_9_1  (
            .in0(N__26168),
            .in1(N__32574),
            .in2(N__29280),
            .in3(N__44570),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_10_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_10_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27008),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_10_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_10_9_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_10_9_3  (
            .in0(N__26511),
            .in1(N__44569),
            .in2(N__33390),
            .in3(N__29331),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44199),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_10_9_5  (
            .in0(N__26682),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_10_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_10_9_6 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_10_9_6  (
            .in0(N__28937),
            .in1(N__32681),
            .in2(N__44596),
            .in3(N__29112),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_10_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_10_9_7 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_10_9_7  (
            .in0(N__32486),
            .in1(N__37877),
            .in2(N__29235),
            .in3(N__44574),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_10_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_10_10_0 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_10_10_0  (
            .in0(N__29364),
            .in1(N__26415),
            .in2(N__29343),
            .in3(N__44531),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_10_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_10_10_1 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_10_10_1  (
            .in0(N__31995),
            .in1(N__26361),
            .in2(N__44584),
            .in3(N__29469),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_10_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_10_10_2 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_10_10_2  (
            .in0(N__29520),
            .in1(N__31899),
            .in2(N__29496),
            .in3(N__44522),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_10_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_10_10_3 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_10_10_3  (
            .in0(N__26298),
            .in1(N__32541),
            .in2(N__44583),
            .in3(N__29253),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_10_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_10_10_4 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_10_10_4  (
            .in0(N__37926),
            .in1(N__28997),
            .in2(N__29481),
            .in3(N__44524),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_10_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_10_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_10_10_5  (
            .in0(N__44518),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_10_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_10_10_6 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_10_10_6  (
            .in0(N__29868),
            .in1(N__32168),
            .in2(N__29532),
            .in3(N__44523),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_10_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_10_10_7 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_10_10_7  (
            .in0(N__32326),
            .in1(N__29433),
            .in2(N__44585),
            .in3(N__29406),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_10_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_10_11_0 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_10_11_0  (
            .in0(N__31847),
            .in1(N__29610),
            .in2(N__44592),
            .in3(N__29583),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_10_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_10_11_1 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_10_11_1  (
            .in0(N__26897),
            .in1(N__44555),
            .in2(N__32208),
            .in3(N__29619),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_10_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_10_11_2 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_10_11_2  (
            .in0(N__29397),
            .in1(N__32270),
            .in2(N__44591),
            .in3(N__29373),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_10_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_10_11_3 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_10_11_3  (
            .in0(N__44928),
            .in1(N__44559),
            .in2(N__40074),
            .in3(N__29559),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_10_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_10_11_4 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_10_11_4  (
            .in0(N__40446),
            .in1(N__26568),
            .in2(N__44593),
            .in3(N__29571),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41697),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_10_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_10_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26896),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_10_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_10_11_7 .LUT_INIT=16'b0011110011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_10_11_7  (
            .in0(N__26846),
            .in1(N__29664),
            .in2(N__29637),
            .in3(N__44554),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_10_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_10_12_0 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_10_12_0  (
            .in0(N__26728),
            .in1(N__44587),
            .in2(N__29307),
            .in3(N__33443),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26727),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_12_2 .LUT_INIT=16'b0000000111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_10_12_2  (
            .in0(N__27345),
            .in1(N__27500),
            .in2(N__27197),
            .in3(N__26769),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49193),
            .ce(),
            .sr(N__48441));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_10_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_10_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_10_12_3 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_10_12_3  (
            .in0(N__27497),
            .in1(N__27347),
            .in2(N__26712),
            .in3(N__27188),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49193),
            .ce(),
            .sr(N__48441));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_10_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_10_12_4 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_10_12_4  (
            .in0(N__27343),
            .in1(N__27498),
            .in2(N__27195),
            .in3(N__26703),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49193),
            .ce(),
            .sr(N__48441));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_12_6 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_10_12_6  (
            .in0(N__27344),
            .in1(N__27499),
            .in2(N__27196),
            .in3(N__26697),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49193),
            .ce(),
            .sr(N__48441));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_10_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_10_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_10_12_7 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_10_12_7  (
            .in0(N__27496),
            .in1(N__27346),
            .in2(N__27213),
            .in3(N__27187),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49193),
            .ce(),
            .sr(N__48441));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_10_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_10_13_0 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_10_13_0  (
            .in0(N__28025),
            .in1(N__26939),
            .in2(N__27978),
            .in3(N__27687),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_13_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_10_13_2  (
            .in0(N__27743),
            .in1(N__26930),
            .in2(N__30066),
            .in3(N__26976),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_13_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_10_13_3  (
            .in0(N__26958),
            .in1(N__30082),
            .in2(N__26964),
            .in3(N__31376),
            .lcout(\phase_controller_inst1.stoper_hc.N_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_10_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_10_13_4 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_10_13_4  (
            .in0(N__26948),
            .in1(N__26940),
            .in2(N__30690),
            .in3(N__31112),
            .lcout(elapsed_time_ns_1_RNIJEKEE1_0_2),
            .ltout(elapsed_time_ns_1_RNIJEKEE1_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_10_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_10_13_5 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26961),
            .in3(N__30149),
            .lcout(\phase_controller_inst1.stoper_hc.N_284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_13_6 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_10_13_6  (
            .in0(N__30150),
            .in1(N__30083),
            .in2(N__26952),
            .in3(N__29687),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_10_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_10_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_10_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_10_13_7  (
            .in0(N__28005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49185),
            .ce(N__28623),
            .sr(N__48453));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_14_0 .LUT_INIT=16'b0011001110111011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_10_14_0  (
            .in0(N__30323),
            .in1(N__27744),
            .in2(_gnd_net_),
            .in3(N__26931),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_10_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_10_14_1 .LUT_INIT=16'b0000000011011100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_10_14_1  (
            .in0(N__30062),
            .in1(N__27627),
            .in2(N__27603),
            .in3(N__31346),
            .lcout(\phase_controller_inst1.stoper_hc.N_326 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_10_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_10_14_2 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__30189),
            .in2(N__27600),
            .in3(N__33183),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_10_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_10_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_10_14_3 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_10_14_3  (
            .in0(N__30190),
            .in1(N__33306),
            .in2(N__27588),
            .in3(N__27581),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49177),
            .ce(N__34502),
            .sr(N__48460));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_10_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_10_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_10_14_7 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_10_14_7  (
            .in0(N__33184),
            .in1(N__33307),
            .in2(N__33034),
            .in3(N__27570),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49177),
            .ce(N__34502),
            .sr(N__48460));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_10_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_10_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_10_15_0  (
            .in0(N__29924),
            .in1(N__28760),
            .in2(N__28812),
            .in3(N__30296),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_10_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_10_15_1 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_10_15_1  (
            .in0(N__31099),
            .in1(N__27540),
            .in2(N__30685),
            .in3(N__28811),
            .lcout(elapsed_time_ns_1_RNIAMU8E1_0_27),
            .ltout(elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_15_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_10_15_2  (
            .in0(N__30362),
            .in1(N__27794),
            .in2(N__27534),
            .in3(N__27674),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_10_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_10_15_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_10_15_3  (
            .in0(N__30677),
            .in1(N__30114),
            .in2(N__31122),
            .in3(N__29721),
            .lcout(elapsed_time_ns_1_RNIOJKEE1_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_10_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_10_15_4 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_10_15_4  (
            .in0(N__31103),
            .in1(N__27531),
            .in2(N__30686),
            .in3(N__30870),
            .lcout(elapsed_time_ns_1_RNI6IU8E1_0_23),
            .ltout(elapsed_time_ns_1_RNI6IU8E1_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_15_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27699),
            .in3(N__27806),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_10_15_6  (
            .in0(N__27641),
            .in1(N__30453),
            .in2(N__27696),
            .in3(N__27693),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_10_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_10_15_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_10_15_7  (
            .in0(N__27860),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27917),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_10_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_10_16_0 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_10_16_0  (
            .in0(N__30852),
            .in1(N__30663),
            .in2(N__27678),
            .in3(N__31066),
            .lcout(elapsed_time_ns_1_RNI9LU8E1_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_10_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_10_16_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_10_16_1  (
            .in0(N__27705),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30253),
            .lcout(elapsed_time_ns_1_RNIDDC6P1_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_10_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_10_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_10_16_2  (
            .in0(N__29700),
            .in1(N__30696),
            .in2(N__27663),
            .in3(N__27651),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_10_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_10_16_3 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_10_16_3  (
            .in0(N__28637),
            .in1(N__49968),
            .in2(N__27645),
            .in3(N__42450),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_10_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_10_16_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_10_16_4  (
            .in0(N__27642),
            .in1(N__30665),
            .in2(N__31749),
            .in3(N__31068),
            .lcout(elapsed_time_ns_1_RNI5HU8E1_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_10_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_10_16_5 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_10_16_5  (
            .in0(N__30666),
            .in1(N__30058),
            .in2(N__31108),
            .in3(N__30720),
            .lcout(elapsed_time_ns_1_RNI7IT8E1_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_10_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_10_16_6 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_10_16_6  (
            .in0(N__27807),
            .in1(N__30664),
            .in2(N__30888),
            .in3(N__31067),
            .lcout(elapsed_time_ns_1_RNI7JU8E1_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_10_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_10_16_7 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_10_16_7  (
            .in0(N__30662),
            .in1(N__28761),
            .in2(N__31107),
            .in3(N__27795),
            .lcout(elapsed_time_ns_1_RNIBNU8E1_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_10_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_10_17_0 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_10_17_0  (
            .in0(N__28082),
            .in1(N__30667),
            .in2(N__27918),
            .in3(N__31072),
            .lcout(elapsed_time_ns_1_RNIMHKEE1_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_10_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_10_17_1 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_10_17_1  (
            .in0(N__30668),
            .in1(N__31537),
            .in2(N__31109),
            .in3(N__31203),
            .lcout(elapsed_time_ns_1_RNI5GT8E1_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_10_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_10_17_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_10_17_2  (
            .in0(N__30915),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30232),
            .lcout(elapsed_time_ns_1_RNIIIC6P1_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_10_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_10_17_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(N__47630),
            .in2(_gnd_net_),
            .in3(N__27779),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_365_clk ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_365_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_10_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_10_17_4 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_10_17_4  (
            .in0(N__30494),
            .in1(N__31173),
            .in2(N__27783),
            .in3(N__30669),
            .lcout(elapsed_time_ns_1_RNI4FT8E1_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_10_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_10_17_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_10_17_5  (
            .in0(N__48587),
            .in1(N__47631),
            .in2(_gnd_net_),
            .in3(N__27780),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_10_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_10_17_6 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_10_17_6  (
            .in0(N__30468),
            .in1(N__30825),
            .in2(N__27765),
            .in3(N__31073),
            .lcout(elapsed_time_ns_1_RNI4GU8E1_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_10_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_10_17_7 .LUT_INIT=16'b1111111011001110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_10_17_7  (
            .in0(N__27742),
            .in1(N__47632),
            .in2(N__31110),
            .in3(N__31188),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_10_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_10_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_10_18_5 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_10_18_5  (
            .in0(N__28078),
            .in1(N__33310),
            .in2(N__33042),
            .in3(N__33117),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49150),
            .ce(N__34506),
            .sr(N__48492));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_10_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_10_18_6 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_10_18_6  (
            .in0(N__28638),
            .in1(N__30673),
            .in2(N__33180),
            .in3(N__31092),
            .lcout(elapsed_time_ns_1_RNI5IV8E1_0_31),
            .ltout(elapsed_time_ns_1_RNI5IV8E1_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_10_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_10_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_10_18_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_10_18_7  (
            .in0(N__33040),
            .in1(_gnd_net_),
            .in2(N__28056),
            .in3(N__30118),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49150),
            .ce(N__34506),
            .sr(N__48492));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__28049),
            .in2(N__27948),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49144),
            .ce(N__28622),
            .sr(N__48504));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__28001),
            .in2(N__27893),
            .in3(N__27951),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49144),
            .ce(N__28622),
            .sr(N__48504));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__27947),
            .in2(N__27839),
            .in3(N__27897),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49144),
            .ce(N__28622),
            .sr(N__48504));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__28343),
            .in2(N__27894),
            .in3(N__27843),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49144),
            .ce(N__28622),
            .sr(N__48504));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__28316),
            .in2(N__27840),
            .in3(N__27810),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49144),
            .ce(N__28622),
            .sr(N__48504));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__28292),
            .in2(N__28347),
            .in3(N__28320),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49144),
            .ce(N__28622),
            .sr(N__48504));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__28317),
            .in2(N__28268),
            .in3(N__28296),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49144),
            .ce(N__28622),
            .sr(N__48504));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__28293),
            .in2(N__28232),
            .in3(N__28272),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49144),
            .ce(N__28622),
            .sr(N__48504));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__28196),
            .in2(N__28269),
            .in3(N__28239),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49139),
            .ce(N__28621),
            .sr(N__48512));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__28163),
            .in2(N__28236),
            .in3(N__28203),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49139),
            .ce(N__28621),
            .sr(N__48512));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__28136),
            .in2(N__28200),
            .in3(N__28167),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49139),
            .ce(N__28621),
            .sr(N__48512));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__28164),
            .in2(N__28112),
            .in3(N__28140),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49139),
            .ce(N__28621),
            .sr(N__48512));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__28137),
            .in2(N__28586),
            .in3(N__28116),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49139),
            .ce(N__28621),
            .sr(N__48512));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__28550),
            .in2(N__28113),
            .in3(N__28086),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49139),
            .ce(N__28621),
            .sr(N__48512));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__28514),
            .in2(N__28587),
            .in3(N__28557),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49139),
            .ce(N__28621),
            .sr(N__48512));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(N__28487),
            .in2(N__28554),
            .in3(N__28521),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49139),
            .ce(N__28621),
            .sr(N__48512));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__28460),
            .in2(N__28518),
            .in3(N__28491),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49134),
            .ce(N__28619),
            .sr(N__48519));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__28488),
            .in2(N__28436),
            .in3(N__28464),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49134),
            .ce(N__28619),
            .sr(N__48519));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__28461),
            .in2(N__28406),
            .in3(N__28440),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49134),
            .ce(N__28619),
            .sr(N__48519));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__28373),
            .in2(N__28437),
            .in3(N__28410),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49134),
            .ce(N__28619),
            .sr(N__48519));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__28889),
            .in2(N__28407),
            .in3(N__28380),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49134),
            .ce(N__28619),
            .sr(N__48519));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__28865),
            .in2(N__28377),
            .in3(N__28350),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49134),
            .ce(N__28619),
            .sr(N__48519));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__28890),
            .in2(N__28841),
            .in3(N__28869),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49134),
            .ce(N__28619),
            .sr(N__48519));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__28866),
            .in2(N__28793),
            .in3(N__28845),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49134),
            .ce(N__28619),
            .sr(N__48519));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__28736),
            .in2(N__28842),
            .in3(N__28797),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49127),
            .ce(N__28618),
            .sr(N__48525));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__28670),
            .in2(N__28794),
            .in3(N__28740),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49127),
            .ce(N__28618),
            .sr(N__48525));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__28737),
            .in2(N__28716),
            .in3(N__28695),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49127),
            .ce(N__28618),
            .sr(N__48525));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__28692),
            .in2(N__28674),
            .in3(N__28644),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49127),
            .ce(N__28618),
            .sr(N__48525));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28641),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49127),
            .ce(N__28618),
            .sr(N__48525));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_10_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_10_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_10_23_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_10_23_0  (
            .in0(N__33187),
            .in1(N__31431),
            .in2(_gnd_net_),
            .in3(N__31305),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49122),
            .ce(N__32879),
            .sr(N__48530));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_10_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_10_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_10_23_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_10_23_2  (
            .in0(N__33186),
            .in1(N__29083),
            .in2(_gnd_net_),
            .in3(N__31432),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49122),
            .ce(N__32879),
            .sr(N__48530));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_10_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_10_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_10_23_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_10_23_4  (
            .in0(N__33188),
            .in1(N__31489),
            .in2(N__30570),
            .in3(N__31433),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49122),
            .ce(N__32879),
            .sr(N__48530));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_10_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_10_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_10_23_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_10_23_5  (
            .in0(N__31430),
            .in1(N__33189),
            .in2(_gnd_net_),
            .in3(N__30950),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49122),
            .ce(N__32879),
            .sr(N__48530));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_10_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_10_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_10_23_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_10_23_7  (
            .in0(N__31236),
            .in1(N__33190),
            .in2(_gnd_net_),
            .in3(N__33018),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49122),
            .ce(N__32879),
            .sr(N__48530));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_11_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_11_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_11_6_5  (
            .in0(N__29515),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44581),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_11_6_7  (
            .in0(N__29428),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44582),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_7_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__44514),
            .in2(_gnd_net_),
            .in3(N__29362),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28998),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_11_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_11_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28933),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29214),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__29154),
            .in2(_gnd_net_),
            .in3(N__36836),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__29148),
            .in2(_gnd_net_),
            .in3(N__32453),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__29142),
            .in2(_gnd_net_),
            .in3(N__32429),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__29136),
            .in2(_gnd_net_),
            .in3(N__32408),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__29130),
            .in2(_gnd_net_),
            .in3(N__29118),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__32040),
            .in2(_gnd_net_),
            .in3(N__29115),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__32514),
            .in2(_gnd_net_),
            .in3(N__29106),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__31788),
            .in2(_gnd_net_),
            .in3(N__29094),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33402),
            .in3(N__29325),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_8 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__33327),
            .in2(_gnd_net_),
            .in3(N__29310),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__33420),
            .in2(_gnd_net_),
            .in3(N__29295),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__32046),
            .in2(_gnd_net_),
            .in3(N__29283),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_11_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_11_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__32052),
            .in2(_gnd_net_),
            .in3(N__29268),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_11_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_11_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__29265),
            .in2(_gnd_net_),
            .in3(N__29247),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__32503),
            .in2(_gnd_net_),
            .in3(N__29238),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__32479),
            .in2(_gnd_net_),
            .in3(N__29226),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__29867),
            .in2(_gnd_net_),
            .in3(N__29523),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__29516),
            .in2(_gnd_net_),
            .in3(N__29484),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__37922),
            .in2(_gnd_net_),
            .in3(N__29472),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__31994),
            .in2(_gnd_net_),
            .in3(N__29463),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__29460),
            .in2(_gnd_net_),
            .in3(N__29436),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__29429),
            .in2(_gnd_net_),
            .in3(N__29400),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__29396),
            .in2(_gnd_net_),
            .in3(N__29367),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__29363),
            .in2(_gnd_net_),
            .in3(N__29334),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__29663),
            .in2(_gnd_net_),
            .in3(N__29622),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32204),
            .in3(N__29613),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__29609),
            .in2(_gnd_net_),
            .in3(N__29577),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__29825),
            .in2(_gnd_net_),
            .in3(N__29574),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__40445),
            .in2(_gnd_net_),
            .in3(N__29565),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__44282),
            .in2(_gnd_net_),
            .in3(N__29562),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__44924),
            .in2(_gnd_net_),
            .in3(N__29553),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_11_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_11_11_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_11_11_7  (
            .in0(N__31971),
            .in1(N__44400),
            .in2(_gnd_net_),
            .in3(N__29550),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_12_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_12_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_11_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29901),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49186),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_12_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_12_1  (
            .in0(N__44380),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_11_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_11_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_11_12_2  (
            .in0(N__29866),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44374),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_11_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_11_12_3 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_11_12_3  (
            .in0(N__44740),
            .in1(N__44283),
            .in2(N__44474),
            .in3(N__29844),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_11_12_5  (
            .in0(N__44375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29826),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_11_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_11_12_6 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_11_12_6  (
            .in0(N__29804),
            .in1(N__44376),
            .in2(N__29763),
            .in3(N__29760),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_11_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_11_13_5 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_11_13_5  (
            .in0(N__33291),
            .in1(N__33185),
            .in2(N__33019),
            .in3(N__32930),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49178),
            .ce(N__34574),
            .sr(N__48442));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_11_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_11_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_11_14_0  (
            .in0(N__29742),
            .in1(N__29720),
            .in2(N__30810),
            .in3(N__30350),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_11_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_11_14_3 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_11_14_3  (
            .in0(N__31345),
            .in1(N__33181),
            .in2(N__30087),
            .in3(N__29688),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_11_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_11_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_11_14_4 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_11_14_4  (
            .in0(N__30162),
            .in1(N__32999),
            .in2(N__30129),
            .in3(N__33308),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49169),
            .ce(N__34558),
            .sr(N__48454));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_11_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_11_14_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_11_14_5  (
            .in0(N__31231),
            .in1(N__30122),
            .in2(N__30006),
            .in3(N__30322),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_11_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_11_14_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_11_14_6  (
            .in0(N__30063),
            .in1(_gnd_net_),
            .in2(N__30009),
            .in3(N__31344),
            .lcout(\phase_controller_inst1.stoper_hc.N_328 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_11_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_11_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_11_14_7 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_11_14_7  (
            .in0(N__30005),
            .in1(N__32998),
            .in2(N__29985),
            .in3(N__33182),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49169),
            .ce(N__34558),
            .sr(N__48454));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__30389),
            .in2(_gnd_net_),
            .in3(N__30407),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_15_2 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_15_2  (
            .in0(N__34441),
            .in1(N__30408),
            .in2(N__33792),
            .in3(N__30390),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49161),
            .ce(),
            .sr(N__48461));
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_11_15_4 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_11_15_4  (
            .in0(N__30443),
            .in1(N__33800),
            .in2(N__29981),
            .in3(N__30391),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49161),
            .ce(),
            .sr(N__48461));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_11_15_6 .LUT_INIT=16'b1011000010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_11_15_6  (
            .in0(N__29950),
            .in1(N__33801),
            .in2(N__30447),
            .in3(N__30392),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49161),
            .ce(),
            .sr(N__48461));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_11_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_11_16_0 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_11_16_0  (
            .in0(N__29928),
            .in1(N__30657),
            .in2(N__31104),
            .in3(N__29907),
            .lcout(elapsed_time_ns_1_RNICOU8E1_0_29),
            .ltout(elapsed_time_ns_1_RNICOU8E1_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_11_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_11_16_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_11_16_1  (
            .in0(N__30278),
            .in1(N__30467),
            .in2(N__30456),
            .in3(N__30581),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_11_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_11_16_2 .LUT_INIT=16'b1111111101110101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_11_16_2  (
            .in0(N__30442),
            .in1(N__35142),
            .in2(N__33819),
            .in3(N__35171),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_11_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_11_16_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30399),
            .in3(N__30396),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_11_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_11_16_4 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_11_16_4  (
            .in0(N__31056),
            .in1(N__30906),
            .in2(N__30366),
            .in3(N__30661),
            .lcout(elapsed_time_ns_1_RNI8KU8E1_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_11_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_11_16_5 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_11_16_5  (
            .in0(N__30656),
            .in1(N__31055),
            .in2(N__30562),
            .in3(N__30351),
            .lcout(elapsed_time_ns_1_RNI2DT8E1_0_10),
            .ltout(elapsed_time_ns_1_RNI2DT8E1_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_11_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_11_16_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_11_16_6  (
            .in0(N__30489),
            .in1(N__31524),
            .in2(N__30333),
            .in3(N__30522),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_11_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_11_16_7 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_11_16_7  (
            .in0(N__30279),
            .in1(N__30300),
            .in2(N__30684),
            .in3(N__31057),
            .lcout(elapsed_time_ns_1_RNI4HV8E1_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_11_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_11_17_0 .LUT_INIT=16'b1011101111111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_11_17_0  (
            .in0(N__47677),
            .in1(N__30270),
            .in2(N__30194),
            .in3(N__31085),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_11_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_11_17_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30258),
            .in3(N__30254),
            .lcout(elapsed_time_ns_1_RNIP93CP1_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_11_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_11_17_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_11_17_2  (
            .in0(N__31155),
            .in1(N__30671),
            .in2(N__30538),
            .in3(N__31081),
            .lcout(elapsed_time_ns_1_RNI3ET8E1_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_11_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_11_17_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_11_17_3  (
            .in0(N__30672),
            .in1(N__31235),
            .in2(N__31111),
            .in3(N__30806),
            .lcout(elapsed_time_ns_1_RNIPKKEE1_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_11_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_11_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_11_17_4  (
            .in0(N__30785),
            .in1(N__30758),
            .in2(N__30744),
            .in3(N__30716),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_11_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_11_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_11_17_5  (
            .in0(N__31731),
            .in1(N__30834),
            .in2(N__30699),
            .in3(N__31140),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_11_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_11_17_6 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_11_17_6  (
            .in0(N__30582),
            .in1(N__30670),
            .in2(N__31782),
            .in3(N__31080),
            .lcout(elapsed_time_ns_1_RNI3FU8E1_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_11_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_11_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_11_18_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_11_18_0  (
            .in0(N__33225),
            .in1(N__30566),
            .in2(N__31505),
            .in3(N__31398),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49145),
            .ce(N__34559),
            .sr(N__48480));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_11_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_11_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_11_18_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_11_18_1  (
            .in0(N__31395),
            .in1(N__31502),
            .in2(N__30540),
            .in3(N__33228),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49145),
            .ce(N__34559),
            .sr(N__48480));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_11_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_11_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_11_18_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_11_18_2  (
            .in0(N__33226),
            .in1(N__30493),
            .in2(N__31506),
            .in3(N__31399),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49145),
            .ce(N__34559),
            .sr(N__48480));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_11_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_11_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_11_18_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_11_18_3  (
            .in0(N__31396),
            .in1(N__33227),
            .in2(N__31542),
            .in3(N__31503),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49145),
            .ce(N__34559),
            .sr(N__48480));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_11_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_11_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_11_18_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_11_18_4  (
            .in0(N__33223),
            .in1(N__31397),
            .in2(_gnd_net_),
            .in3(N__31304),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49145),
            .ce(N__34559),
            .sr(N__48480));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_18_5 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_11_18_5  (
            .in0(N__34216),
            .in1(N__31268),
            .in2(N__34254),
            .in3(N__31254),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_11_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_11_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_11_18_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_11_18_6  (
            .in0(N__33224),
            .in1(N__33036),
            .in2(_gnd_net_),
            .in3(N__31230),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49145),
            .ce(N__34559),
            .sr(N__48480));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_11_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_11_19_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_11_19_3  (
            .in0(N__31199),
            .in1(N__31184),
            .in2(N__31172),
            .in3(N__31151),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_11_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_11_19_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_11_19_7  (
            .in0(N__46885),
            .in1(N__42129),
            .in2(_gnd_net_),
            .in3(N__46320),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_11_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_11_20_4 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_11_20_4  (
            .in0(N__31760),
            .in1(N__31123),
            .in2(N__30954),
            .in3(N__47700),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_20_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_11_20_5  (
            .in0(N__30899),
            .in1(N__30881),
            .in2(N__30869),
            .in3(N__30845),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_11_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_11_20_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_11_20_6  (
            .in0(N__30821),
            .in1(N__31772),
            .in2(N__31761),
            .in3(N__31742),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_21_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_11_21_4  (
            .in0(N__35557),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34357),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_1_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(N__35615),
            .in2(_gnd_net_),
            .in3(N__31613),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(N__34309),
            .in2(_gnd_net_),
            .in3(N__31567),
            .lcout(\phase_controller_inst1.start_timer_hc_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_11_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_11_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_11_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31644),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49123),
            .ce(),
            .sr(N__48520));
    defparam \phase_controller_inst1.state_3_LC_11_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_11_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_11_22_5 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst1.state_3_LC_11_22_5  (
            .in0(N__35628),
            .in1(N__35424),
            .in2(N__31620),
            .in3(N__31682),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49123),
            .ce(),
            .sr(N__48520));
    defparam \phase_controller_inst1.start_timer_hc_LC_11_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_11_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_11_22_6 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_11_22_6  (
            .in0(N__35408),
            .in1(N__31662),
            .in2(N__31650),
            .in3(N__31656),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49123),
            .ce(),
            .sr(N__48520));
    defparam \phase_controller_inst1.state_2_LC_11_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_11_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_11_23_6 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst1.state_2_LC_11_23_6  (
            .in0(N__31612),
            .in1(N__34302),
            .in2(N__31578),
            .in3(N__35629),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49118),
            .ce(),
            .sr(N__48526));
    defparam \phase_controller_inst1.state_1_LC_11_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_11_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_11_24_5 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \phase_controller_inst1.state_1_LC_11_24_5  (
            .in0(N__31577),
            .in1(N__34308),
            .in2(N__35568),
            .in3(N__34361),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49115),
            .ce(),
            .sr(N__48531));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32034),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__40922),
            .in2(_gnd_net_),
            .in3(N__37507),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_395_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_12_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_6_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37545),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32004),
            .ce(),
            .sr(N__48396));
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_6_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_12_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37546),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32004),
            .ce(),
            .sr(N__48396));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_12_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_12_7_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(N__44513),
            .in2(_gnd_net_),
            .in3(N__31987),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_12_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_12_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31968),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31900),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_12_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_12_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31843),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_8_1  (
            .in0(N__32650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_12_8_2  (
            .in0(N__32327),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_12_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_12_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_12_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32265),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_12_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_12_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43579),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_6  (
            .in0(N__32197),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44495),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32163),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_9_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_9_0  (
            .in0(N__44512),
            .in1(N__32108),
            .in2(N__32351),
            .in3(N__32073),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32566),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32599),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32344),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32669),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_12_9_5  (
            .in0(N__32507),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44510),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_12_9_6  (
            .in0(N__44511),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32487),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_10_0  (
            .in0(N__34686),
            .in1(N__32466),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__34680),
            .in2(_gnd_net_),
            .in3(N__32439),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__49192),
            .ce(),
            .sr(N__48413));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__34671),
            .in2(_gnd_net_),
            .in3(N__32415),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__49192),
            .ce(),
            .sr(N__48413));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__34767),
            .in2(_gnd_net_),
            .in3(N__32391),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__49192),
            .ce(),
            .sr(N__48413));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__34758),
            .in2(_gnd_net_),
            .in3(N__32361),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__49192),
            .ce(),
            .sr(N__48413));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__34749),
            .in2(_gnd_net_),
            .in3(N__32331),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__49192),
            .ce(),
            .sr(N__48413));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(N__34740),
            .in2(_gnd_net_),
            .in3(N__32658),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__49192),
            .ce(),
            .sr(N__48413));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__34731),
            .in2(_gnd_net_),
            .in3(N__32625),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__49192),
            .ce(),
            .sr(N__48413));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__34722),
            .in2(_gnd_net_),
            .in3(N__32622),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__49184),
            .ce(),
            .sr(N__48418));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__34713),
            .in2(_gnd_net_),
            .in3(N__32619),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__49184),
            .ce(),
            .sr(N__48418));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__34704),
            .in2(_gnd_net_),
            .in3(N__32616),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__49184),
            .ce(),
            .sr(N__48418));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__34812),
            .in2(_gnd_net_),
            .in3(N__32577),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__49184),
            .ce(),
            .sr(N__48418));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__34803),
            .in2(_gnd_net_),
            .in3(N__32544),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__49184),
            .ce(),
            .sr(N__48418));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_12_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_12_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_12_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__33408),
            .in2(_gnd_net_),
            .in3(N__32520),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__49184),
            .ce(),
            .sr(N__48418));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_12_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_12_11_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__34791),
            .in2(_gnd_net_),
            .in3(N__32517),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49184),
            .ce(),
            .sr(N__48418));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33431),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_12_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__37290),
            .in2(_gnd_net_),
            .in3(N__37314),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__37242),
            .in2(_gnd_net_),
            .in3(N__37266),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34790),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33379),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_12_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_12_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_12_12_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_12_12_5  (
            .in0(N__33380),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49176),
            .ce(),
            .sr(N__48426));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(N__33340),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_12_13_1  (
            .in0(N__33292),
            .in1(N__33243),
            .in2(N__33041),
            .in3(N__32934),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49168),
            .ce(N__32899),
            .sr(N__48431));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__33603),
            .in2(N__33594),
            .in3(N__33784),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__33585),
            .in2(N__33579),
            .in3(N__33999),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__33570),
            .in2(N__33564),
            .in3(N__33974),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__33555),
            .in2(N__33546),
            .in3(N__33954),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__33537),
            .in2(N__33522),
            .in3(N__33936),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_12_14_5  (
            .in0(N__33918),
            .in1(N__33504),
            .in2(N__33513),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__33498),
            .in2(N__33483),
            .in3(N__33900),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__33471),
            .in2(N__33459),
            .in3(N__33882),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__33768),
            .in2(N__33756),
            .in3(N__33861),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__33747),
            .in2(N__33738),
            .in3(N__34173),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__33717),
            .in2(N__33729),
            .in3(N__34155),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__33711),
            .in2(N__33702),
            .in3(N__34137),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__33681),
            .in2(N__33693),
            .in3(N__34119),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_12_15_5  (
            .in0(N__34101),
            .in1(N__33675),
            .in2(N__33660),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__33651),
            .in2(N__33639),
            .in3(N__34083),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__33630),
            .in2(N__33618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__33840),
            .in2(N__33831),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__35463),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__35286),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35253),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35217),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__35181),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__35172),
            .in2(N__35118),
            .in3(N__33807),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33804),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__33791),
            .in2(N__34011),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_12_17_1  (
            .in0(N__34551),
            .in1(N__33998),
            .in2(_gnd_net_),
            .in3(N__33984),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49143),
            .ce(),
            .sr(N__48467));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_17_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_12_17_2  (
            .in0(N__34555),
            .in1(N__33981),
            .in2(N__33975),
            .in3(N__33957),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49143),
            .ce(),
            .sr(N__48467));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_12_17_3  (
            .in0(N__34552),
            .in1(N__33953),
            .in2(_gnd_net_),
            .in3(N__33939),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49143),
            .ce(),
            .sr(N__48467));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_12_17_4  (
            .in0(N__34556),
            .in1(N__33935),
            .in2(_gnd_net_),
            .in3(N__33921),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49143),
            .ce(),
            .sr(N__48467));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_12_17_5  (
            .in0(N__34553),
            .in1(N__33917),
            .in2(_gnd_net_),
            .in3(N__33903),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49143),
            .ce(),
            .sr(N__48467));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_12_17_6  (
            .in0(N__34557),
            .in1(N__33899),
            .in2(_gnd_net_),
            .in3(N__33885),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49143),
            .ce(),
            .sr(N__48467));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_12_17_7  (
            .in0(N__34554),
            .in1(N__33878),
            .in2(_gnd_net_),
            .in3(N__33864),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49143),
            .ce(),
            .sr(N__48467));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_12_18_0  (
            .in0(N__34531),
            .in1(N__33857),
            .in2(_gnd_net_),
            .in3(N__33843),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49138),
            .ce(),
            .sr(N__48473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_12_18_1  (
            .in0(N__34508),
            .in1(N__34172),
            .in2(_gnd_net_),
            .in3(N__34158),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49138),
            .ce(),
            .sr(N__48473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_12_18_2  (
            .in0(N__34528),
            .in1(N__34154),
            .in2(_gnd_net_),
            .in3(N__34140),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49138),
            .ce(),
            .sr(N__48473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_12_18_3  (
            .in0(N__34509),
            .in1(N__34136),
            .in2(_gnd_net_),
            .in3(N__34122),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49138),
            .ce(),
            .sr(N__48473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_12_18_4  (
            .in0(N__34529),
            .in1(N__34118),
            .in2(_gnd_net_),
            .in3(N__34104),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49138),
            .ce(),
            .sr(N__48473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_12_18_5  (
            .in0(N__34510),
            .in1(N__34100),
            .in2(_gnd_net_),
            .in3(N__34086),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49138),
            .ce(),
            .sr(N__48473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_12_18_6  (
            .in0(N__34530),
            .in1(N__34082),
            .in2(_gnd_net_),
            .in3(N__34068),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49138),
            .ce(),
            .sr(N__48473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_12_18_7  (
            .in0(N__34511),
            .in1(N__34055),
            .in2(_gnd_net_),
            .in3(N__34041),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49138),
            .ce(),
            .sr(N__48473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_12_19_0  (
            .in0(N__34512),
            .in1(N__34028),
            .in2(_gnd_net_),
            .in3(N__34014),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49133),
            .ce(),
            .sr(N__48481));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_12_19_1  (
            .in0(N__34567),
            .in1(N__34246),
            .in2(_gnd_net_),
            .in3(N__34227),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49133),
            .ce(),
            .sr(N__48481));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_12_19_2  (
            .in0(N__34513),
            .in1(N__34217),
            .in2(_gnd_net_),
            .in3(N__34197),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49133),
            .ce(),
            .sr(N__48481));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_12_19_3  (
            .in0(N__34568),
            .in1(N__35475),
            .in2(_gnd_net_),
            .in3(N__34194),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49133),
            .ce(),
            .sr(N__48481));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_12_19_4  (
            .in0(N__34514),
            .in1(N__35487),
            .in2(_gnd_net_),
            .in3(N__34191),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49133),
            .ce(),
            .sr(N__48481));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_12_19_5  (
            .in0(N__34569),
            .in1(N__35298),
            .in2(_gnd_net_),
            .in3(N__34188),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49133),
            .ce(),
            .sr(N__48481));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_12_19_6  (
            .in0(N__34515),
            .in1(N__35310),
            .in2(_gnd_net_),
            .in3(N__34185),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49133),
            .ce(),
            .sr(N__48481));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_12_19_7  (
            .in0(N__34570),
            .in1(N__35277),
            .in2(_gnd_net_),
            .in3(N__34182),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49133),
            .ce(),
            .sr(N__48481));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_12_20_0  (
            .in0(N__34560),
            .in1(N__35265),
            .in2(_gnd_net_),
            .in3(N__34179),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49126),
            .ce(),
            .sr(N__48493));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_12_20_1  (
            .in0(N__34571),
            .in1(N__35241),
            .in2(_gnd_net_),
            .in3(N__34176),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49126),
            .ce(),
            .sr(N__48493));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_12_20_2  (
            .in0(N__34561),
            .in1(N__35229),
            .in2(_gnd_net_),
            .in3(N__34587),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49126),
            .ce(),
            .sr(N__48493));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_12_20_3  (
            .in0(N__34572),
            .in1(N__35193),
            .in2(_gnd_net_),
            .in3(N__34584),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49126),
            .ce(),
            .sr(N__48493));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_12_20_4  (
            .in0(N__34562),
            .in1(N__35205),
            .in2(_gnd_net_),
            .in3(N__34581),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49126),
            .ce(),
            .sr(N__48493));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_12_20_5  (
            .in0(N__34573),
            .in1(N__35138),
            .in2(_gnd_net_),
            .in3(N__34578),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49126),
            .ce(),
            .sr(N__48493));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_12_20_6  (
            .in0(N__34563),
            .in1(N__35164),
            .in2(_gnd_net_),
            .in3(N__34368),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49126),
            .ce(),
            .sr(N__48493));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(N__35668),
            .in2(_gnd_net_),
            .in3(N__35449),
            .lcout(\phase_controller_inst1.time_passed_RNI7NN7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_0_LC_12_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_12_22_0 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \phase_controller_inst1.state_0_LC_12_22_0  (
            .in0(N__35450),
            .in1(N__34365),
            .in2(N__35571),
            .in3(N__35669),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49117),
            .ce(),
            .sr(N__48513));
    defparam \phase_controller_inst1.T12_LC_12_26_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.T12_LC_12_26_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T12_LC_12_26_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst1.T12_LC_12_26_3  (
            .in0(N__34322),
            .in1(N__34311),
            .in2(_gnd_net_),
            .in3(N__35564),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48535));
    defparam \phase_controller_inst1.T01_LC_12_26_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_12_26_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_12_26_5 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \phase_controller_inst1.T01_LC_12_26_5  (
            .in0(N__35645),
            .in1(N__34310),
            .in2(_gnd_net_),
            .in3(N__34265),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49110),
            .ce(),
            .sr(N__48535));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_5_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_13_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35813),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_6_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_6_1  (
            .in0(N__35757),
            .in1(N__35814),
            .in2(_gnd_net_),
            .in3(N__35784),
            .lcout(\current_shift_inst.timer_s1.N_167_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_7_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_7_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__40734),
            .in2(N__36020),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49216),
            .ce(N__44133),
            .sr(N__48397));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_7_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__44159),
            .in2(N__35994),
            .in3(N__34605),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49216),
            .ce(N__44133),
            .sr(N__48397));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_7_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__35960),
            .in2(N__36021),
            .in3(N__34602),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49216),
            .ce(N__44133),
            .sr(N__48397));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_7_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__35990),
            .in2(N__35939),
            .in3(N__34599),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49216),
            .ce(N__44133),
            .sr(N__48397));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_7_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_7_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__35961),
            .in2(N__35912),
            .in3(N__34596),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49216),
            .ce(N__44133),
            .sr(N__48397));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_7_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_7_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__35882),
            .in2(N__35940),
            .in3(N__34593),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49216),
            .ce(N__44133),
            .sr(N__48397));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_7_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_7_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(N__35845),
            .in2(N__35913),
            .in3(N__34590),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49216),
            .ce(N__44133),
            .sr(N__48397));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_7_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_7_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__36226),
            .in2(N__35883),
            .in3(N__34632),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49216),
            .ce(N__44133),
            .sr(N__48397));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(N__36206),
            .in2(N__35853),
            .in3(N__34629),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49208),
            .ce(N__44131),
            .sr(N__48400));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__36182),
            .in2(N__36237),
            .in3(N__34626),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49208),
            .ce(N__44131),
            .sr(N__48400));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__36207),
            .in2(N__36161),
            .in3(N__34623),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49208),
            .ce(N__44131),
            .sr(N__48400));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__36183),
            .in2(N__36131),
            .in3(N__34620),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49208),
            .ce(N__44131),
            .sr(N__48400));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(N__36104),
            .in2(N__36162),
            .in3(N__34617),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49208),
            .ce(N__44131),
            .sr(N__48400));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__36080),
            .in2(N__36132),
            .in3(N__34614),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49208),
            .ce(N__44131),
            .sr(N__48400));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__36105),
            .in2(N__36050),
            .in3(N__34611),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49208),
            .ce(N__44131),
            .sr(N__48400));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__36469),
            .in2(N__36084),
            .in3(N__34608),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49208),
            .ce(N__44131),
            .sr(N__48400));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__36449),
            .in2(N__36054),
            .in3(N__34662),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49203),
            .ce(N__44130),
            .sr(N__48403));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__36425),
            .in2(N__36480),
            .in3(N__34659),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49203),
            .ce(N__44130),
            .sr(N__48403));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__36450),
            .in2(N__36404),
            .in3(N__34656),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49203),
            .ce(N__44130),
            .sr(N__48403));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__36426),
            .in2(N__36374),
            .in3(N__34653),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49203),
            .ce(N__44130),
            .sr(N__48403));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__36347),
            .in2(N__36405),
            .in3(N__34650),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49203),
            .ce(N__44130),
            .sr(N__48403));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__36326),
            .in2(N__36375),
            .in3(N__34647),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49203),
            .ce(N__44130),
            .sr(N__48403));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__36348),
            .in2(N__36293),
            .in3(N__34644),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49203),
            .ce(N__44130),
            .sr(N__48403));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__36256),
            .in2(N__36327),
            .in3(N__34641),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49203),
            .ce(N__44130),
            .sr(N__48403));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__36297),
            .in2(N__36737),
            .in3(N__34638),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49197),
            .ce(N__44128),
            .sr(N__48405));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__36710),
            .in2(N__36267),
            .in3(N__34635),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49197),
            .ce(N__44128),
            .sr(N__48405));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__36690),
            .in2(N__36738),
            .in3(N__34695),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49197),
            .ce(N__44128),
            .sr(N__48405));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__36711),
            .in2(N__36546),
            .in3(N__34692),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49197),
            .ce(N__44128),
            .sr(N__48405));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34689),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40204),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40397),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_13_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_13_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39851),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_13_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_13_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__36744),
            .in2(N__36791),
            .in3(N__36787),
            .lcout(\current_shift_inst.control_input_18 ),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_11_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__36804),
            .in2(_gnd_net_),
            .in3(N__34674),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_11_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__36768),
            .in2(_gnd_net_),
            .in3(N__34665),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_11_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__36762),
            .in2(_gnd_net_),
            .in3(N__34761),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_11_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__36756),
            .in2(_gnd_net_),
            .in3(N__34752),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_11_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__36750),
            .in2(_gnd_net_),
            .in3(N__34743),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_11_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__36954),
            .in2(_gnd_net_),
            .in3(N__34734),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_11_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__36948),
            .in2(_gnd_net_),
            .in3(N__34725),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_12_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__36939),
            .in2(_gnd_net_),
            .in3(N__34716),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_12_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__36930),
            .in2(_gnd_net_),
            .in3(N__34707),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__36924),
            .in2(_gnd_net_),
            .in3(N__34698),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_12_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__38451),
            .in2(_gnd_net_),
            .in3(N__34806),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__36798),
            .in2(_gnd_net_),
            .in3(N__34797),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_13_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_13_12_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__38529),
            .in2(_gnd_net_),
            .in3(N__34794),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_13_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_13_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_13_13_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_13_13_7  (
            .in0(N__40868),
            .in1(N__49596),
            .in2(N__42339),
            .in3(N__46823),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49179),
            .ce(N__48802),
            .sr(N__48427));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(N__34889),
            .in2(_gnd_net_),
            .in3(N__34868),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_13_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_13_14_1 .LUT_INIT=16'b1111011111110101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_13_14_1  (
            .in0(N__34917),
            .in1(N__37458),
            .in2(N__37491),
            .in3(N__35337),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_13_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_13_14_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34779),
            .in3(N__34890),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_LC_13_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_13_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_13_14_4 .LUT_INIT=16'b1000101011111010;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_13_14_4  (
            .in0(N__34776),
            .in1(N__35322),
            .in2(N__34898),
            .in3(N__34919),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49170),
            .ce(),
            .sr(N__48432));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_14_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_14_5  (
            .in0(N__34916),
            .in1(N__34775),
            .in2(_gnd_net_),
            .in3(N__34964),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_6 .LUT_INIT=16'b1011101000001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_13_14_6  (
            .in0(N__34984),
            .in1(N__35321),
            .in2(N__34899),
            .in3(N__34918),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49170),
            .ce(),
            .sr(N__48432));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_13_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_13_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_13_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34965),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49170),
            .ce(),
            .sr(N__48432));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_13_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_13_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_13_15_0 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_13_15_0  (
            .in0(N__34891),
            .in1(N__34869),
            .in2(N__36918),
            .in3(N__50170),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49162),
            .ce(),
            .sr(N__48443));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_13_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_13_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_13_15_5 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_13_15_5  (
            .in0(N__40914),
            .in1(N__37563),
            .in2(_gnd_net_),
            .in3(N__37523),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49162),
            .ce(),
            .sr(N__48443));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__47490),
            .in2(N__34857),
            .in3(N__36913),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__50436),
            .in2(N__34848),
            .in3(N__36888),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_16_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_16_2  (
            .in0(N__36861),
            .in1(N__46503),
            .in2(N__34839),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__50295),
            .in2(N__34830),
            .in3(N__37119),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(N__46518),
            .in2(N__34821),
            .in3(N__37101),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_16_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_16_5  (
            .in0(N__37083),
            .in1(N__35061),
            .in2(N__46668),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(N__47502),
            .in2(N__35055),
            .in3(N__37065),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_16_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_16_7  (
            .in0(N__37047),
            .in1(N__45021),
            .in2(N__35046),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_17_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_17_0  (
            .in0(N__37029),
            .in1(N__38700),
            .in2(N__35037),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__37380),
            .in2(N__35028),
            .in3(N__37011),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_17_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_17_2  (
            .in0(N__36990),
            .in1(N__38745),
            .in2(N__35019),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__38733),
            .in2(N__35010),
            .in3(N__36972),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__38439),
            .in2(N__34998),
            .in3(N__37218),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_17_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_17_5  (
            .in0(N__37200),
            .in1(N__37371),
            .in2(N__35100),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__35091),
            .in2(N__37395),
            .in3(N__37182),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__38829),
            .in2(N__38769),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__38688),
            .in2(N__38625),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__35106),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35496),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__37401),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__35085),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__35073),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__37483),
            .in2(N__37437),
            .in3(N__35328),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35325),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_19_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__35309),
            .in2(_gnd_net_),
            .in3(N__35297),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_19_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_13_19_1  (
            .in0(N__35276),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35264),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_13_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_13_19_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_13_19_2  (
            .in0(N__35240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35228),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_19_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__35204),
            .in2(_gnd_net_),
            .in3(N__35192),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_19_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__35163),
            .in2(_gnd_net_),
            .in3(N__35137),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_13_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_13_19_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__37134),
            .in2(_gnd_net_),
            .in3(N__37152),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_13_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_13_19_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_13_19_6  (
            .in0(N__37356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37338),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_13_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_13_20_0 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_13_20_0  (
            .in0(N__37652),
            .in1(N__37607),
            .in2(_gnd_net_),
            .in3(N__35352),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_20_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_13_20_1  (
            .in0(N__35353),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37653),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_20_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_13_20_2  (
            .in0(N__37737),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37719),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_20_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__35486),
            .in2(_gnd_net_),
            .in3(N__35474),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_21_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_21_0 .LUT_INIT=16'b1101000011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_13_21_0  (
            .in0(N__39456),
            .in1(N__35451),
            .in2(N__37659),
            .in3(N__37631),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49128),
            .ce(),
            .sr(N__48494));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35355),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49128),
            .ce(),
            .sr(N__48494));
    defparam \phase_controller_inst1.start_timer_tr_LC_13_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_21_3 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_13_21_3  (
            .in0(N__35433),
            .in1(N__35423),
            .in2(N__35412),
            .in3(N__35354),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49128),
            .ce(),
            .sr(N__48494));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_13_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_13_22_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(N__37751),
            .in2(_gnd_net_),
            .in3(N__37766),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_22_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(N__37818),
            .in2(_gnd_net_),
            .in3(N__37832),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_22_7  (
            .in0(N__35800),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35775),
            .lcout(\current_shift_inst.timer_s1.N_166_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_LC_13_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_23_0 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_23_0  (
            .in0(N__35779),
            .in1(N__35750),
            .in2(_gnd_net_),
            .in3(N__35806),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49119),
            .ce(),
            .sr(N__48514));
    defparam \current_shift_inst.stop_timer_s1_LC_13_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_13_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_13_23_1 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_13_23_1  (
            .in0(N__35749),
            .in1(N__35780),
            .in2(N__35652),
            .in3(N__35723),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49119),
            .ce(),
            .sr(N__48514));
    defparam \current_shift_inst.start_timer_s1_LC_13_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_13_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_13_24_2 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_13_24_2  (
            .in0(N__35716),
            .in1(N__35748),
            .in2(_gnd_net_),
            .in3(N__35651),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49116),
            .ce(),
            .sr(N__48521));
    defparam \phase_controller_inst1.S1_LC_13_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_13_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35650),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49114),
            .ce(),
            .sr(N__48527));
    defparam \phase_controller_inst1.T23_LC_13_26_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.T23_LC_13_26_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T23_LC_13_26_0 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst1.T23_LC_13_26_0  (
            .in0(N__35690),
            .in1(N__35569),
            .in2(_gnd_net_),
            .in3(N__35678),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49113),
            .ce(),
            .sr(N__48532));
    defparam \phase_controller_inst1.T45_LC_13_26_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.T45_LC_13_26_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T45_LC_13_26_3 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \phase_controller_inst1.T45_LC_13_26_3  (
            .in0(N__35679),
            .in1(N__35582),
            .in2(_gnd_net_),
            .in3(N__35649),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49113),
            .ce(),
            .sr(N__48532));
    defparam \phase_controller_inst1.S2_LC_13_27_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_27_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_27_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_27_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35570),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49111),
            .ce(),
            .sr(N__48536));
    defparam \current_shift_inst.timer_s1.counter_0_LC_14_5_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_14_5_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_14_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_14_5_0  (
            .in0(N__36667),
            .in1(N__40726),
            .in2(_gnd_net_),
            .in3(N__35499),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__49232),
            .ce(N__36523),
            .sr(N__48393));
    defparam \current_shift_inst.timer_s1.counter_1_LC_14_5_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_14_5_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_14_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_14_5_1  (
            .in0(N__36629),
            .in1(N__44155),
            .in2(_gnd_net_),
            .in3(N__36024),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__49232),
            .ce(N__36523),
            .sr(N__48393));
    defparam \current_shift_inst.timer_s1.counter_2_LC_14_5_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_14_5_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_14_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_14_5_2  (
            .in0(N__36668),
            .in1(N__36013),
            .in2(_gnd_net_),
            .in3(N__35997),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__49232),
            .ce(N__36523),
            .sr(N__48393));
    defparam \current_shift_inst.timer_s1.counter_3_LC_14_5_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_14_5_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_14_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_14_5_3  (
            .in0(N__36630),
            .in1(N__35986),
            .in2(_gnd_net_),
            .in3(N__35964),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__49232),
            .ce(N__36523),
            .sr(N__48393));
    defparam \current_shift_inst.timer_s1.counter_4_LC_14_5_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_14_5_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_14_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_14_5_4  (
            .in0(N__36669),
            .in1(N__35959),
            .in2(_gnd_net_),
            .in3(N__35943),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__49232),
            .ce(N__36523),
            .sr(N__48393));
    defparam \current_shift_inst.timer_s1.counter_5_LC_14_5_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_14_5_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_14_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_14_5_5  (
            .in0(N__36631),
            .in1(N__35932),
            .in2(_gnd_net_),
            .in3(N__35916),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__49232),
            .ce(N__36523),
            .sr(N__48393));
    defparam \current_shift_inst.timer_s1.counter_6_LC_14_5_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_14_5_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_14_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_14_5_6  (
            .in0(N__36670),
            .in1(N__35900),
            .in2(_gnd_net_),
            .in3(N__35886),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__49232),
            .ce(N__36523),
            .sr(N__48393));
    defparam \current_shift_inst.timer_s1.counter_7_LC_14_5_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_14_5_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_14_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_14_5_7  (
            .in0(N__36632),
            .in1(N__35875),
            .in2(_gnd_net_),
            .in3(N__35856),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__49232),
            .ce(N__36523),
            .sr(N__48393));
    defparam \current_shift_inst.timer_s1.counter_8_LC_14_6_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_14_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_14_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_14_6_0  (
            .in0(N__36666),
            .in1(N__35849),
            .in2(_gnd_net_),
            .in3(N__35829),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__49227),
            .ce(N__36524),
            .sr(N__48394));
    defparam \current_shift_inst.timer_s1.counter_9_LC_14_6_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_14_6_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_14_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_14_6_1  (
            .in0(N__36636),
            .in1(N__36230),
            .in2(_gnd_net_),
            .in3(N__36210),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__49227),
            .ce(N__36524),
            .sr(N__48394));
    defparam \current_shift_inst.timer_s1.counter_10_LC_14_6_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_14_6_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_14_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_14_6_2  (
            .in0(N__36663),
            .in1(N__36200),
            .in2(_gnd_net_),
            .in3(N__36186),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__49227),
            .ce(N__36524),
            .sr(N__48394));
    defparam \current_shift_inst.timer_s1.counter_11_LC_14_6_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_14_6_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_14_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_14_6_3  (
            .in0(N__36633),
            .in1(N__36181),
            .in2(_gnd_net_),
            .in3(N__36165),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__49227),
            .ce(N__36524),
            .sr(N__48394));
    defparam \current_shift_inst.timer_s1.counter_12_LC_14_6_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_14_6_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_14_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_14_6_4  (
            .in0(N__36664),
            .in1(N__36149),
            .in2(_gnd_net_),
            .in3(N__36135),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__49227),
            .ce(N__36524),
            .sr(N__48394));
    defparam \current_shift_inst.timer_s1.counter_13_LC_14_6_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_14_6_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_14_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_14_6_5  (
            .in0(N__36634),
            .in1(N__36124),
            .in2(_gnd_net_),
            .in3(N__36108),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__49227),
            .ce(N__36524),
            .sr(N__48394));
    defparam \current_shift_inst.timer_s1.counter_14_LC_14_6_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_14_6_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_14_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_14_6_6  (
            .in0(N__36665),
            .in1(N__36103),
            .in2(_gnd_net_),
            .in3(N__36087),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__49227),
            .ce(N__36524),
            .sr(N__48394));
    defparam \current_shift_inst.timer_s1.counter_15_LC_14_6_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_14_6_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_14_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_14_6_7  (
            .in0(N__36635),
            .in1(N__36073),
            .in2(_gnd_net_),
            .in3(N__36057),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__49227),
            .ce(N__36524),
            .sr(N__48394));
    defparam \current_shift_inst.timer_s1.counter_16_LC_14_7_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_14_7_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_14_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_14_7_0  (
            .in0(N__36646),
            .in1(N__36049),
            .in2(_gnd_net_),
            .in3(N__36027),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__49221),
            .ce(N__36516),
            .sr(N__48395));
    defparam \current_shift_inst.timer_s1.counter_17_LC_14_7_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_14_7_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_14_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_14_7_1  (
            .in0(N__36654),
            .in1(N__36473),
            .in2(_gnd_net_),
            .in3(N__36453),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__49221),
            .ce(N__36516),
            .sr(N__48395));
    defparam \current_shift_inst.timer_s1.counter_18_LC_14_7_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_14_7_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_14_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_14_7_2  (
            .in0(N__36647),
            .in1(N__36443),
            .in2(_gnd_net_),
            .in3(N__36429),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__49221),
            .ce(N__36516),
            .sr(N__48395));
    defparam \current_shift_inst.timer_s1.counter_19_LC_14_7_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_14_7_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_14_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_14_7_3  (
            .in0(N__36655),
            .in1(N__36424),
            .in2(_gnd_net_),
            .in3(N__36408),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__49221),
            .ce(N__36516),
            .sr(N__48395));
    defparam \current_shift_inst.timer_s1.counter_20_LC_14_7_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_14_7_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_14_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_14_7_4  (
            .in0(N__36648),
            .in1(N__36392),
            .in2(_gnd_net_),
            .in3(N__36378),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__49221),
            .ce(N__36516),
            .sr(N__48395));
    defparam \current_shift_inst.timer_s1.counter_21_LC_14_7_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_14_7_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_14_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_14_7_5  (
            .in0(N__36656),
            .in1(N__36367),
            .in2(_gnd_net_),
            .in3(N__36351),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__49221),
            .ce(N__36516),
            .sr(N__48395));
    defparam \current_shift_inst.timer_s1.counter_22_LC_14_7_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_14_7_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_14_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_14_7_6  (
            .in0(N__36649),
            .in1(N__36346),
            .in2(_gnd_net_),
            .in3(N__36330),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__49221),
            .ce(N__36516),
            .sr(N__48395));
    defparam \current_shift_inst.timer_s1.counter_23_LC_14_7_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_14_7_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_14_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_14_7_7  (
            .in0(N__36657),
            .in1(N__36319),
            .in2(_gnd_net_),
            .in3(N__36300),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__49221),
            .ce(N__36516),
            .sr(N__48395));
    defparam \current_shift_inst.timer_s1.counter_24_LC_14_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_14_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_14_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_14_8_0  (
            .in0(N__36650),
            .in1(N__36292),
            .in2(_gnd_net_),
            .in3(N__36270),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__49217),
            .ce(N__36528),
            .sr(N__48398));
    defparam \current_shift_inst.timer_s1.counter_25_LC_14_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_14_8_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_14_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_14_8_1  (
            .in0(N__36671),
            .in1(N__36260),
            .in2(_gnd_net_),
            .in3(N__36240),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__49217),
            .ce(N__36528),
            .sr(N__48398));
    defparam \current_shift_inst.timer_s1.counter_26_LC_14_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_14_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_14_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_14_8_2  (
            .in0(N__36651),
            .in1(N__36730),
            .in2(_gnd_net_),
            .in3(N__36714),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__49217),
            .ce(N__36528),
            .sr(N__48398));
    defparam \current_shift_inst.timer_s1.counter_27_LC_14_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_14_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_14_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_14_8_3  (
            .in0(N__36672),
            .in1(N__36709),
            .in2(_gnd_net_),
            .in3(N__36693),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__49217),
            .ce(N__36528),
            .sr(N__48398));
    defparam \current_shift_inst.timer_s1.counter_28_LC_14_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_14_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_14_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_14_8_4  (
            .in0(N__36652),
            .in1(N__36689),
            .in2(_gnd_net_),
            .in3(N__36675),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__49217),
            .ce(N__36528),
            .sr(N__48398));
    defparam \current_shift_inst.timer_s1.counter_29_LC_14_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_14_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_14_8_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_14_8_5  (
            .in0(N__36542),
            .in1(N__36653),
            .in2(_gnd_net_),
            .in3(N__36549),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49217),
            .ce(N__36528),
            .sr(N__48398));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_9_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_14_9_0  (
            .in0(N__39791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44652),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_14_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_14_9_2 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_14_9_2  (
            .in0(N__44052),
            .in1(N__41064),
            .in2(_gnd_net_),
            .in3(N__40666),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_9_3  (
            .in0(N__38162),
            .in1(_gnd_net_),
            .in2(N__36486),
            .in3(N__36813),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_9_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__38163),
            .in2(N__36483),
            .in3(N__41616),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46162),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_9_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_14_9_6  (
            .in0(N__44053),
            .in1(_gnd_net_),
            .in2(N__41761),
            .in3(N__41735),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41752),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_10_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_14_10_0  (
            .in0(N__40244),
            .in1(N__45443),
            .in2(_gnd_net_),
            .in3(N__41473),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40243),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_10_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_14_10_2  (
            .in0(N__43414),
            .in1(N__44036),
            .in2(_gnd_net_),
            .in3(N__43385),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43413),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_10_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_14_10_4  (
            .in0(N__39683),
            .in1(N__44037),
            .in2(_gnd_net_),
            .in3(N__41157),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39682),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_14_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_14_10_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_14_10_6  (
            .in0(N__41886),
            .in1(N__38418),
            .in2(_gnd_net_),
            .in3(N__38494),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_14_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_14_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_14_10_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36843),
            .in3(N__36792),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49204),
            .ce(),
            .sr(N__48404));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39973),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49198),
            .ce(N__44129),
            .sr(N__48406));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_14_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_14_12_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_14_12_0  (
            .in0(N__38403),
            .in1(N__41862),
            .in2(_gnd_net_),
            .in3(N__38496),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38514),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_14_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_14_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38495),
            .lcout(\current_shift_inst.N_1460_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_12_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_14_12_3  (
            .in0(N__38497),
            .in1(N__38391),
            .in2(_gnd_net_),
            .in3(N__42063),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_14_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_14_12_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_14_12_4  (
            .in0(N__38379),
            .in1(N__42048),
            .in2(_gnd_net_),
            .in3(N__38498),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_12_5 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_12_5  (
            .in0(N__38367),
            .in1(N__38512),
            .in2(_gnd_net_),
            .in3(N__42021),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_12_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_12_6  (
            .in0(N__38513),
            .in1(N__42000),
            .in2(_gnd_net_),
            .in3(N__38601),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_12_7 .LUT_INIT=16'b0010011100100111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_14_12_7  (
            .in0(N__38499),
            .in1(N__38589),
            .in2(N__41976),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_13_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_14_13_0  (
            .in0(N__41946),
            .in1(N__38577),
            .in2(_gnd_net_),
            .in3(N__38518),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_13_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_14_13_1  (
            .in0(N__38519),
            .in1(N__41916),
            .in2(_gnd_net_),
            .in3(N__38565),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_13_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_14_13_2  (
            .in0(N__41901),
            .in1(N__38553),
            .in2(_gnd_net_),
            .in3(N__38520),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_14_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_14_13_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_14_13_3  (
            .in0(N__38521),
            .in1(N__42300),
            .in2(_gnd_net_),
            .in3(N__38541),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__36914),
            .in2(N__36897),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_14_1  (
            .in0(N__50260),
            .in1(N__36887),
            .in2(_gnd_net_),
            .in3(N__36873),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49180),
            .ce(),
            .sr(N__48428));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_14_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_14_2  (
            .in0(N__50277),
            .in1(N__36860),
            .in2(N__36870),
            .in3(N__36846),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49180),
            .ce(),
            .sr(N__48428));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_14_3  (
            .in0(N__50261),
            .in1(N__37118),
            .in2(_gnd_net_),
            .in3(N__37104),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49180),
            .ce(),
            .sr(N__48428));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_14_4  (
            .in0(N__50278),
            .in1(N__37100),
            .in2(_gnd_net_),
            .in3(N__37086),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49180),
            .ce(),
            .sr(N__48428));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_14_5  (
            .in0(N__50262),
            .in1(N__37082),
            .in2(_gnd_net_),
            .in3(N__37068),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49180),
            .ce(),
            .sr(N__48428));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_14_6  (
            .in0(N__50279),
            .in1(N__37064),
            .in2(_gnd_net_),
            .in3(N__37050),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49180),
            .ce(),
            .sr(N__48428));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_14_7  (
            .in0(N__50263),
            .in1(N__37046),
            .in2(_gnd_net_),
            .in3(N__37032),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49180),
            .ce(),
            .sr(N__48428));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_15_0  (
            .in0(N__50163),
            .in1(N__37028),
            .in2(_gnd_net_),
            .in3(N__37014),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49171),
            .ce(),
            .sr(N__48433));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_15_1  (
            .in0(N__50156),
            .in1(N__37007),
            .in2(_gnd_net_),
            .in3(N__36993),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49171),
            .ce(),
            .sr(N__48433));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_15_2  (
            .in0(N__50160),
            .in1(N__36989),
            .in2(_gnd_net_),
            .in3(N__36975),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49171),
            .ce(),
            .sr(N__48433));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_15_3  (
            .in0(N__50157),
            .in1(N__36971),
            .in2(_gnd_net_),
            .in3(N__36957),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49171),
            .ce(),
            .sr(N__48433));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_15_4  (
            .in0(N__50161),
            .in1(N__37217),
            .in2(_gnd_net_),
            .in3(N__37203),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49171),
            .ce(),
            .sr(N__48433));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_15_5  (
            .in0(N__50158),
            .in1(N__37199),
            .in2(_gnd_net_),
            .in3(N__37185),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49171),
            .ce(),
            .sr(N__48433));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_15_6  (
            .in0(N__50162),
            .in1(N__37181),
            .in2(_gnd_net_),
            .in3(N__37167),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49171),
            .ce(),
            .sr(N__48433));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_15_7  (
            .in0(N__50159),
            .in1(N__38812),
            .in2(_gnd_net_),
            .in3(N__37164),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49171),
            .ce(),
            .sr(N__48433));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_16_0  (
            .in0(N__50237),
            .in1(N__38784),
            .in2(_gnd_net_),
            .in3(N__37161),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49163),
            .ce(),
            .sr(N__48444));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_16_1  (
            .in0(N__50245),
            .in1(N__38660),
            .in2(_gnd_net_),
            .in3(N__37158),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49163),
            .ce(),
            .sr(N__48444));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_16_2  (
            .in0(N__50238),
            .in1(N__38643),
            .in2(_gnd_net_),
            .in3(N__37155),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49163),
            .ce(),
            .sr(N__48444));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_16_3  (
            .in0(N__50246),
            .in1(N__37151),
            .in2(_gnd_net_),
            .in3(N__37137),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49163),
            .ce(),
            .sr(N__48444));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_16_4  (
            .in0(N__50239),
            .in1(N__37133),
            .in2(_gnd_net_),
            .in3(N__37359),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49163),
            .ce(),
            .sr(N__48444));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_16_5  (
            .in0(N__50247),
            .in1(N__37355),
            .in2(_gnd_net_),
            .in3(N__37341),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49163),
            .ce(),
            .sr(N__48444));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_16_6  (
            .in0(N__50240),
            .in1(N__37337),
            .in2(_gnd_net_),
            .in3(N__37323),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49163),
            .ce(),
            .sr(N__48444));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_16_7  (
            .in0(N__50248),
            .in1(N__37427),
            .in2(_gnd_net_),
            .in3(N__37320),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49163),
            .ce(),
            .sr(N__48444));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_17_0  (
            .in0(N__50241),
            .in1(N__37413),
            .in2(_gnd_net_),
            .in3(N__37317),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49156),
            .ce(),
            .sr(N__48455));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_17_1  (
            .in0(N__50249),
            .in1(N__37307),
            .in2(_gnd_net_),
            .in3(N__37293),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49156),
            .ce(),
            .sr(N__48455));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_17_2  (
            .in0(N__50242),
            .in1(N__37283),
            .in2(_gnd_net_),
            .in3(N__37269),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49156),
            .ce(),
            .sr(N__48455));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_17_3  (
            .in0(N__50250),
            .in1(N__37259),
            .in2(_gnd_net_),
            .in3(N__37245),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49156),
            .ce(),
            .sr(N__48455));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_17_4  (
            .in0(N__50243),
            .in1(N__37235),
            .in2(_gnd_net_),
            .in3(N__37221),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49156),
            .ce(),
            .sr(N__48455));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_17_5  (
            .in0(N__50251),
            .in1(N__37457),
            .in2(_gnd_net_),
            .in3(N__37569),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49156),
            .ce(),
            .sr(N__48455));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_17_6  (
            .in0(N__50244),
            .in1(N__37484),
            .in2(_gnd_net_),
            .in3(N__37566),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49156),
            .ce(),
            .sr(N__48455));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_18_0 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_14_18_0  (
            .in0(N__37559),
            .in1(N__40921),
            .in2(_gnd_net_),
            .in3(N__37527),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_396_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_14_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_14_18_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_14_18_2  (
            .in0(N__37482),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37456),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_18_6 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_18_6  (
            .in0(N__37428),
            .in1(N__37412),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_14_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_14_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_14_19_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_14_19_0  (
            .in0(N__42404),
            .in1(N__49566),
            .in2(N__46890),
            .in3(N__46817),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49146),
            .ce(N__50259),
            .sr(N__48468));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_14_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_14_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_14_19_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_14_19_2  (
            .in0(N__40866),
            .in1(N__49564),
            .in2(N__42266),
            .in3(N__46815),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49146),
            .ce(N__50259),
            .sr(N__48468));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_14_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_14_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_14_19_6 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_14_19_6  (
            .in0(N__40867),
            .in1(N__49565),
            .in2(N__42180),
            .in3(N__46816),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49146),
            .ce(N__50259),
            .sr(N__48468));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_14_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_14_20_0 .LUT_INIT=16'b1100111011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_14_20_0  (
            .in0(N__39471),
            .in1(N__39359),
            .in2(N__39330),
            .in3(N__37654),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_20_1 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__37625),
            .in2(N__37671),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_14_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_14_20_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_14_20_2  (
            .in0(N__37626),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37667),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_20_3 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_14_20_3  (
            .in0(N__37668),
            .in1(N__37630),
            .in2(N__38957),
            .in3(N__48666),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49140),
            .ce(),
            .sr(N__48474));
    defparam \phase_controller_inst1.stoper_tr.running_LC_14_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_14_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_14_20_4 .LUT_INIT=16'b1011111100110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_14_20_4  (
            .in0(N__39455),
            .in1(N__37655),
            .in2(N__37632),
            .in3(N__37608),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49140),
            .ce(),
            .sr(N__48474));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__37596),
            .in2(N__38958),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_14_21_1  (
            .in0(N__48667),
            .in1(N__38922),
            .in2(_gnd_net_),
            .in3(N__37590),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49135),
            .ce(),
            .sr(N__48482));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_21_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_14_21_2  (
            .in0(N__48753),
            .in1(N__38901),
            .in2(N__37587),
            .in3(N__37578),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49135),
            .ce(),
            .sr(N__48482));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_14_21_3  (
            .in0(N__48668),
            .in1(N__38880),
            .in2(_gnd_net_),
            .in3(N__37575),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49135),
            .ce(),
            .sr(N__48482));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_14_21_4  (
            .in0(N__48754),
            .in1(N__38859),
            .in2(_gnd_net_),
            .in3(N__37572),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49135),
            .ce(),
            .sr(N__48482));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_14_21_5  (
            .in0(N__48669),
            .in1(N__39167),
            .in2(_gnd_net_),
            .in3(N__37698),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49135),
            .ce(),
            .sr(N__48482));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_14_21_6  (
            .in0(N__48755),
            .in1(N__39135),
            .in2(_gnd_net_),
            .in3(N__37695),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49135),
            .ce(),
            .sr(N__48482));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_21_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_14_21_7  (
            .in0(N__48670),
            .in1(N__39117),
            .in2(_gnd_net_),
            .in3(N__37692),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49135),
            .ce(),
            .sr(N__48482));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_22_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_14_22_0  (
            .in0(N__48763),
            .in1(N__39090),
            .in2(_gnd_net_),
            .in3(N__37689),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49129),
            .ce(),
            .sr(N__48495));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_14_22_1  (
            .in0(N__48749),
            .in1(N__39069),
            .in2(_gnd_net_),
            .in3(N__37686),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49129),
            .ce(),
            .sr(N__48495));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_14_22_2  (
            .in0(N__48760),
            .in1(N__39021),
            .in2(_gnd_net_),
            .in3(N__37683),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49129),
            .ce(),
            .sr(N__48495));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_14_22_3  (
            .in0(N__48750),
            .in1(N__39000),
            .in2(_gnd_net_),
            .in3(N__37680),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49129),
            .ce(),
            .sr(N__48495));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_14_22_4  (
            .in0(N__48761),
            .in1(N__38979),
            .in2(_gnd_net_),
            .in3(N__37677),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49129),
            .ce(),
            .sr(N__48495));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_14_22_5  (
            .in0(N__48751),
            .in1(N__39249),
            .in2(_gnd_net_),
            .in3(N__37674),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49129),
            .ce(),
            .sr(N__48495));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_14_22_6  (
            .in0(N__48762),
            .in1(N__39216),
            .in2(_gnd_net_),
            .in3(N__37782),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49129),
            .ce(),
            .sr(N__48495));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_14_22_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_14_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_14_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_14_22_7  (
            .in0(N__48752),
            .in1(N__39424),
            .in2(_gnd_net_),
            .in3(N__37779),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49129),
            .ce(),
            .sr(N__48495));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_14_23_0  (
            .in0(N__48745),
            .in1(N__39408),
            .in2(_gnd_net_),
            .in3(N__37776),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49124),
            .ce(),
            .sr(N__48505));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_14_23_1  (
            .in0(N__48812),
            .in1(N__39561),
            .in2(_gnd_net_),
            .in3(N__37773),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49124),
            .ce(),
            .sr(N__48505));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_14_23_2  (
            .in0(N__48746),
            .in1(N__39579),
            .in2(_gnd_net_),
            .in3(N__37770),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49124),
            .ce(),
            .sr(N__48505));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_14_23_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_14_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_14_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_14_23_3  (
            .in0(N__48813),
            .in1(N__37767),
            .in2(_gnd_net_),
            .in3(N__37755),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49124),
            .ce(),
            .sr(N__48505));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_14_23_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_14_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_14_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_14_23_4  (
            .in0(N__48747),
            .in1(N__37752),
            .in2(_gnd_net_),
            .in3(N__37740),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49124),
            .ce(),
            .sr(N__48505));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_14_23_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_14_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_14_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_14_23_5  (
            .in0(N__48814),
            .in1(N__37736),
            .in2(_gnd_net_),
            .in3(N__37722),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49124),
            .ce(),
            .sr(N__48505));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_14_23_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_14_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_14_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_14_23_6  (
            .in0(N__48748),
            .in1(N__37715),
            .in2(_gnd_net_),
            .in3(N__37701),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49124),
            .ce(),
            .sr(N__48505));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_14_23_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_14_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_14_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_14_23_7  (
            .in0(N__48815),
            .in1(N__37833),
            .in2(_gnd_net_),
            .in3(N__37821),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49124),
            .ce(),
            .sr(N__48505));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_14_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_14_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_14_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_14_24_0  (
            .in0(N__48756),
            .in1(N__37817),
            .in2(_gnd_net_),
            .in3(N__37803),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49120),
            .ce(),
            .sr(N__48515));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_14_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_14_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_14_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_14_24_1  (
            .in0(N__48805),
            .in1(N__39612),
            .in2(_gnd_net_),
            .in3(N__37800),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49120),
            .ce(),
            .sr(N__48515));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_14_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_14_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_14_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_14_24_2  (
            .in0(N__48757),
            .in1(N__39600),
            .in2(_gnd_net_),
            .in3(N__37797),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49120),
            .ce(),
            .sr(N__48515));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_14_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_14_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_14_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_14_24_3  (
            .in0(N__48806),
            .in1(N__39279),
            .in2(_gnd_net_),
            .in3(N__37794),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49120),
            .ce(),
            .sr(N__48515));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_14_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_14_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_14_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_14_24_4  (
            .in0(N__48758),
            .in1(N__39291),
            .in2(_gnd_net_),
            .in3(N__37791),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49120),
            .ce(),
            .sr(N__48515));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_14_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_14_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_14_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_14_24_5  (
            .in0(N__48807),
            .in1(N__39323),
            .in2(_gnd_net_),
            .in3(N__37788),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49120),
            .ce(),
            .sr(N__48515));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_14_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_14_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_14_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_14_24_6  (
            .in0(N__48759),
            .in1(N__39358),
            .in2(_gnd_net_),
            .in3(N__37785),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49120),
            .ce(),
            .sr(N__48515));
    defparam CONSTANT_ONE_LUT4_LC_15_5_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_15_5_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_15_5_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_15_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_15_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_15_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_15_6_0  (
            .in0(_gnd_net_),
            .in1(N__37915),
            .in2(_gnd_net_),
            .in3(N__44580),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37895),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_6_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_6_2  (
            .in0(N__45885),
            .in1(N__45421),
            .in2(N__44676),
            .in3(N__44634),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_6_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_6_3  (
            .in0(N__45418),
            .in1(N__45886),
            .in2(N__40950),
            .in3(N__39525),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_6_4 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_6_4  (
            .in0(N__45884),
            .in1(N__45420),
            .in2(N__43740),
            .in3(N__43775),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_6_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_6_5  (
            .in0(N__45419),
            .in1(N__45887),
            .in2(N__41103),
            .in3(N__41208),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43774),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_7_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_15_7_0  (
            .in0(N__43302),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_7_1  (
            .in0(N__41088),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40692),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_7_3 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_7_3  (
            .in0(N__45422),
            .in1(N__41256),
            .in2(N__40702),
            .in3(N__45882),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_7_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_7_4  (
            .in0(N__45883),
            .in1(N__45423),
            .in2(N__43312),
            .in3(N__43334),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40113),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39514),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_7_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_7_7  (
            .in0(N__41089),
            .in1(N__44055),
            .in2(_gnd_net_),
            .in3(N__41204),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__43841),
            .in2(N__37935),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__38057),
            .in2(N__43899),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__39531),
            .in2(N__38138),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__38061),
            .in2(N__39480),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__39495),
            .in2(N__38139),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__38065),
            .in2(N__39489),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(N__37965),
            .in2(N__38140),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__38069),
            .in2(N__37956),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__38082),
            .in2(N__39624),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__37947),
            .in2(N__38144),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__38070),
            .in2(N__39774),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__37941),
            .in2(N__38141),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__38074),
            .in2(N__39654),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__39636),
            .in2(N__38142),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_9_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__38078),
            .in2(N__39645),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_9_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__39630),
            .in2(N__38143),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__38086),
            .in2(N__39723),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__39714),
            .in2(N__38145),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__38090),
            .in2(N__39756),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__39702),
            .in2(N__38146),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__38094),
            .in2(N__39732),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__39780),
            .in2(N__38147),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__38098),
            .in2(N__39765),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__39708),
            .in2(N__38148),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__38149),
            .in2(N__40143),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__38289),
            .in2(N__38192),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__38153),
            .in2(N__40083),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__39993),
            .in2(N__38193),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__38157),
            .in2(N__39840),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__39888),
            .in2(N__38194),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__38161),
            .in2(N__43884),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_11_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__45393),
            .in2(_gnd_net_),
            .in3(N__38328),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__41633),
            .in2(N__39924),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__44086),
            .in2(N__43266),
            .in3(N__43842),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_12_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_15_12_2  (
            .in0(N__43843),
            .in1(N__45583),
            .in2(N__39960),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__40089),
            .in2(N__45748),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__45587),
            .in2(N__38325),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__38313),
            .in2(N__45749),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(N__45591),
            .in2(N__39906),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__38301),
            .in2(N__45750),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__45637),
            .in2(N__38355),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__39696),
            .in2(N__45840),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__45641),
            .in2(N__40329),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__40335),
            .in2(N__45841),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__45645),
            .in2(N__43626),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__40149),
            .in2(N__45842),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__45649),
            .in2(N__39897),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(N__38340),
            .in2(N__45843),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__45719),
            .in2(N__40170),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__40347),
            .in2(N__45900),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__45723),
            .in2(N__40002),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__38427),
            .in2(N__45901),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__45727),
            .in2(N__39747),
            .in3(N__38406),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__39819),
            .in2(N__45902),
            .in3(N__38394),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__45731),
            .in2(N__46215),
            .in3(N__38382),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__40341),
            .in2(N__45903),
            .in3(N__38370),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__45735),
            .in2(N__40179),
            .in3(N__38358),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__40230),
            .in2(N__45904),
            .in3(N__38592),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__45739),
            .in2(N__40188),
            .in3(N__38580),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__40386),
            .in2(N__45905),
            .in3(N__38568),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__45743),
            .in2(N__39882),
            .in3(N__38556),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__40161),
            .in2(N__45906),
            .in3(N__38544),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_15_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_15_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__45747),
            .in2(N__43800),
            .in3(N__38532),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_15_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_15_15_7 .LUT_INIT=16'b1000101101000111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_15_15_7  (
            .in0(N__39831),
            .in1(N__38528),
            .in2(N__42282),
            .in3(N__38454),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_15_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_15_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_15_16_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_15_16_1  (
            .in0(N__49468),
            .in1(N__42203),
            .in2(N__40860),
            .in3(N__46752),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49172),
            .ce(N__50285),
            .sr(N__48434));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_16_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_15_16_2  (
            .in0(N__46878),
            .in1(N__42397),
            .in2(_gnd_net_),
            .in3(N__42170),
            .lcout(\phase_controller_inst1.stoper_tr.N_242 ),
            .ltout(\phase_controller_inst1.stoper_tr.N_242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_15_16_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_15_16_3  (
            .in0(N__49467),
            .in1(N__42334),
            .in2(N__38748),
            .in3(N__46751),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49172),
            .ce(N__50285),
            .sr(N__48434));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_15_16_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_15_16_4  (
            .in0(N__46749),
            .in1(N__42229),
            .in2(N__40859),
            .in3(N__49469),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49172),
            .ce(N__50285),
            .sr(N__48434));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_15_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_15_16_5 .LUT_INIT=16'b1010101011111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_15_16_5  (
            .in0(N__49466),
            .in1(N__38715),
            .in2(N__42489),
            .in3(N__46748),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_15_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_15_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_15_16_6 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_15_16_6  (
            .in0(N__46750),
            .in1(N__40838),
            .in2(N__38703),
            .in3(N__42123),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49172),
            .ce(N__50285),
            .sr(N__48434));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_15_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_15_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_15_17_1 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_15_17_1  (
            .in0(N__47784),
            .in1(_gnd_net_),
            .in2(N__49598),
            .in3(N__46765),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49164),
            .ce(N__50276),
            .sr(N__48445));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_17_2 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_15_17_2  (
            .in0(N__38609),
            .in1(N__38641),
            .in2(N__38676),
            .in3(N__38659),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_17_3 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_17_3  (
            .in0(N__38672),
            .in1(N__38610),
            .in2(N__38661),
            .in3(N__38642),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_15_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_15_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_15_17_4 .LUT_INIT=16'b0011001100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__49567),
            .in2(N__46807),
            .in3(N__42556),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49164),
            .ce(N__50276),
            .sr(N__48445));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_15_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_15_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_15_17_5 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_15_17_5  (
            .in0(N__42517),
            .in1(_gnd_net_),
            .in2(N__49597),
            .in3(N__46764),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49164),
            .ce(N__50276),
            .sr(N__48445));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_17_6 .LUT_INIT=16'b1111011101010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_17_6  (
            .in0(N__38782),
            .in1(N__38814),
            .in2(N__46446),
            .in3(N__38792),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_17_7 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_17_7  (
            .in0(N__38813),
            .in1(N__46445),
            .in2(N__38796),
            .in3(N__38783),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_15_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_15_18_0 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_15_18_0  (
            .in0(N__42560),
            .in1(N__49860),
            .in2(N__47644),
            .in3(N__42948),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_18_5 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_15_18_5  (
            .in0(N__42978),
            .in1(N__42521),
            .in2(N__49887),
            .in3(N__47611),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_15_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_15_18_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__47822),
            .in2(_gnd_net_),
            .in3(N__38754),
            .lcout(elapsed_time_ns_1_RNIQENQL1_0_9),
            .ltout(elapsed_time_ns_1_RNIQENQL1_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_15_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_15_18_7 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_15_18_7  (
            .in0(N__42834),
            .in1(N__49817),
            .in2(N__38757),
            .in3(N__47610),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_19_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_15_19_0  (
            .in0(N__40864),
            .in1(N__49584),
            .in2(N__42267),
            .in3(N__46813),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49151),
            .ce(N__48803),
            .sr(N__48462));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_15_19_2 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__50386),
            .in2(N__47538),
            .in3(N__49583),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49151),
            .ce(N__48803),
            .sr(N__48462));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_19_3 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_15_19_3  (
            .in0(N__49582),
            .in1(N__49382),
            .in2(N__46551),
            .in3(N__50392),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49151),
            .ce(N__48803),
            .sr(N__48462));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_19_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_15_19_4  (
            .in0(N__46886),
            .in1(N__49585),
            .in2(N__42408),
            .in3(N__46814),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49151),
            .ce(N__48803),
            .sr(N__48462));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_15_19_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_15_19_5  (
            .in0(N__49581),
            .in1(N__47886),
            .in2(_gnd_net_),
            .in3(N__50393),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49151),
            .ce(N__48803),
            .sr(N__48462));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_19_7 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_15_19_7  (
            .in0(N__42168),
            .in1(N__46812),
            .in2(N__49599),
            .in3(N__40865),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49151),
            .ce(N__48803),
            .sr(N__48462));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_20_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_20_0  (
            .in0(N__38947),
            .in1(N__49266),
            .in2(N__38931),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__46644),
            .in2(N__38910),
            .in3(N__38921),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__45057),
            .in2(N__38889),
            .in3(N__38900),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__46656),
            .in2(N__38868),
            .in3(N__38879),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_20_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_20_4  (
            .in0(N__38858),
            .in1(N__38847),
            .in2(N__38841),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(N__46617),
            .in2(N__39153),
            .in3(N__39168),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__39123),
            .in2(N__39144),
            .in3(N__39134),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_20_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_20_7  (
            .in0(N__39116),
            .in1(N__39096),
            .in2(N__39105),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_21_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_21_0  (
            .in0(N__39089),
            .in1(N__40359),
            .in2(N__39078),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_21_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_21_1  (
            .in0(N__39068),
            .in1(N__39057),
            .in2(N__39045),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__39036),
            .in2(N__39009),
            .in3(N__39020),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__40785),
            .in2(N__38988),
            .in3(N__38999),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(N__40377),
            .in2(N__38967),
            .in3(N__38978),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_21_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_21_5  (
            .in0(_gnd_net_),
            .in1(N__39258),
            .in2(N__39237),
            .in3(N__39248),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__39204),
            .in2(N__39228),
            .in3(N__39215),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_21_7  (
            .in0(_gnd_net_),
            .in1(N__39435),
            .in2(N__39393),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__39366),
            .in2(N__39543),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__39198),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_22_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(N__39189),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_22_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(N__39177),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_22_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(N__39588),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_22_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__39267),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(N__39360),
            .in2(N__39303),
            .in3(N__39462),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39459),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_23_0 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_23_0  (
            .in0(N__39406),
            .in1(N__40775),
            .in2(N__39378),
            .in3(N__39426),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_23_1 .LUT_INIT=16'b1111011100110001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_15_23_1  (
            .in0(N__39425),
            .in1(N__39407),
            .in2(N__40779),
            .in3(N__39374),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_15_23_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_15_23_3  (
            .in0(N__49580),
            .in1(N__42525),
            .in2(_gnd_net_),
            .in3(N__46824),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49130),
            .ce(N__48804),
            .sr(N__48496));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_15_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_15_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_15_23_5 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_15_23_5  (
            .in0(N__40745),
            .in1(N__39577),
            .in2(N__40766),
            .in3(N__39559),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_15_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_15_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_15_24_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_15_24_2  (
            .in0(_gnd_net_),
            .in1(N__39354),
            .in2(_gnd_net_),
            .in3(N__39322),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_15_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_15_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_15_24_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_15_24_4  (
            .in0(_gnd_net_),
            .in1(N__39290),
            .in2(_gnd_net_),
            .in3(N__39278),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_15_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_15_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_15_24_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_15_24_6  (
            .in0(N__39611),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39599),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_24_7 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_15_24_7  (
            .in0(N__40746),
            .in1(N__39578),
            .in2(N__40767),
            .in3(N__39560),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_6_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_16_6_7  (
            .in0(N__45409),
            .in1(N__45988),
            .in2(N__40130),
            .in3(N__40979),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_7_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_16_7_0  (
            .in0(N__40943),
            .in1(N__45410),
            .in2(N__46013),
            .in3(N__39524),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_7_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_7_1  (
            .in0(N__39941),
            .in1(N__44038),
            .in2(_gnd_net_),
            .in3(N__41009),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39940),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_7_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_7_3  (
            .in0(N__39523),
            .in1(N__44040),
            .in2(_gnd_net_),
            .in3(N__40942),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_7_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_7_4  (
            .in0(N__44041),
            .in1(N__40703),
            .in2(_gnd_net_),
            .in3(N__41251),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_7_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_7_5  (
            .in0(N__40123),
            .in1(N__44039),
            .in2(_gnd_net_),
            .in3(N__40978),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_7_6 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_16_7_6  (
            .in0(N__45986),
            .in1(N__41149),
            .in2(N__39684),
            .in3(N__45411),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_16_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_16_7_7 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_16_7_7  (
            .in0(N__45412),
            .in1(N__39681),
            .in2(N__41156),
            .in3(N__45987),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43488),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_8_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_8_1  (
            .in0(N__44802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_8_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_8_2  (
            .in0(N__43683),
            .in1(N__44047),
            .in2(_gnd_net_),
            .in3(N__43642),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_8_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_16_8_3  (
            .in0(N__44049),
            .in1(N__46095),
            .in2(_gnd_net_),
            .in3(N__46045),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_8_4 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_16_8_4  (
            .in0(N__43456),
            .in1(N__44048),
            .in2(_gnd_net_),
            .in3(N__43489),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_8_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_8_5  (
            .in0(N__44050),
            .in1(N__43773),
            .in2(_gnd_net_),
            .in3(N__43736),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_8_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_8_6  (
            .in0(N__43313),
            .in1(N__44045),
            .in2(_gnd_net_),
            .in3(N__43327),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_8_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_8_7  (
            .in0(N__44046),
            .in1(_gnd_net_),
            .in2(N__44812),
            .in3(N__44773),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_9_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_9_0  (
            .in0(N__44022),
            .in1(_gnd_net_),
            .in2(N__46273),
            .in3(N__46231),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_9_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_9_1  (
            .in0(N__44212),
            .in1(N__44019),
            .in2(_gnd_net_),
            .in3(N__44236),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_9_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_16_9_2  (
            .in0(N__45345),
            .in1(N__45876),
            .in2(N__45122),
            .in3(N__45095),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_9_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_9_3  (
            .in0(N__45094),
            .in1(N__44021),
            .in2(_gnd_net_),
            .in3(N__45115),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_9_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_9_4  (
            .in0(N__44017),
            .in1(N__43607),
            .in2(_gnd_net_),
            .in3(N__43553),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_9_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_9_5  (
            .in0(N__46189),
            .in1(N__44018),
            .in2(_gnd_net_),
            .in3(N__46138),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_9_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_9_6  (
            .in0(N__44023),
            .in1(N__44994),
            .in2(_gnd_net_),
            .in3(N__44956),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_9_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_9_7  (
            .in0(N__44671),
            .in1(N__44020),
            .in2(_gnd_net_),
            .in3(N__44626),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_10_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_10_0  (
            .in0(N__45301),
            .in1(N__39863),
            .in2(N__45974),
            .in3(N__41357),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_10_1 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_10_1  (
            .in0(N__41358),
            .in1(N__45300),
            .in2(N__39864),
            .in3(N__45848),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_10_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_10_2  (
            .in0(N__45299),
            .in1(N__39859),
            .in2(_gnd_net_),
            .in3(N__41356),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_10_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__45302),
            .in2(_gnd_net_),
            .in3(N__45844),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_16_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_16_10_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_16_10_4  (
            .in0(N__45297),
            .in1(N__39806),
            .in2(N__45975),
            .in3(N__41549),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_10_5 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_16_10_5  (
            .in0(N__41550),
            .in1(N__45298),
            .in2(N__39807),
            .in3(N__45852),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_10_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_10_6  (
            .in0(N__44024),
            .in1(N__39802),
            .in2(_gnd_net_),
            .in3(N__41548),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_10_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_10_7  (
            .in0(N__39980),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49218),
            .ce(N__44134),
            .sr(N__48399));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_11_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_16_11_0  (
            .in0(N__45251),
            .in1(N__45672),
            .in2(N__41390),
            .in3(N__40415),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_11_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_11_1  (
            .in0(N__45392),
            .in1(N__40414),
            .in2(_gnd_net_),
            .in3(N__41383),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39987),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49209),
            .ce(N__44132),
            .sr(N__48401));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_16_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_16_11_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_16_11_3  (
            .in0(N__45673),
            .in1(N__45250),
            .in2(N__39951),
            .in3(N__41018),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_11_4 .LUT_INIT=16'b1010001110100011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_16_11_4  (
            .in0(N__41019),
            .in1(N__39947),
            .in2(N__45364),
            .in3(N__45674),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_11_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_11_5 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_16_11_5  (
            .in0(N__39915),
            .in1(N__40668),
            .in2(_gnd_net_),
            .in3(N__45249),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_16_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_16_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41063),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_16_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_16_11_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__45245),
            .in2(N__39909),
            .in3(N__40667),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_12_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_16_12_0  (
            .in0(N__45805),
            .in1(N__45339),
            .in2(N__43428),
            .in3(N__43386),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_12_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_16_12_1  (
            .in0(N__45341),
            .in1(N__45803),
            .in2(N__46112),
            .in3(N__46056),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_12_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_12_2  (
            .in0(N__44900),
            .in1(N__45343),
            .in2(_gnd_net_),
            .in3(N__44858),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_12_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_12_3  (
            .in0(N__45344),
            .in1(N__45801),
            .in2(N__44862),
            .in3(N__44901),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_16_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_16_12_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_16_12_4  (
            .in0(N__45802),
            .in1(N__45340),
            .in2(N__43503),
            .in3(N__43464),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_12_5 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_12_5  (
            .in0(N__41657),
            .in1(N__44051),
            .in2(_gnd_net_),
            .in3(N__41701),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_12_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_16_12_6  (
            .in0(N__45804),
            .in1(N__45338),
            .in2(N__40134),
            .in3(N__40986),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_12_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_12_7  (
            .in0(N__45342),
            .in1(N__40222),
            .in2(_gnd_net_),
            .in3(N__41431),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_16_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_16_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40072),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_13_1 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_16_13_1  (
            .in0(N__40223),
            .in1(N__45679),
            .in2(N__45444),
            .in3(N__41438),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_13_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_16_13_2  (
            .in0(N__40256),
            .in1(N__45399),
            .in2(N__45874),
            .in3(N__41480),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_16_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_16_13_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_16_13_3  (
            .in0(N__45397),
            .in1(N__45685),
            .in2(N__44220),
            .in3(N__44247),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_16_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_16_13_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_16_13_4  (
            .in0(N__46193),
            .in1(N__45396),
            .in2(N__45875),
            .in3(N__46146),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_13_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_16_13_5  (
            .in0(N__45398),
            .in1(N__45675),
            .in2(N__45006),
            .in3(N__44964),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_16_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_16_13_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_16_13_6  (
            .in0(N__45681),
            .in1(N__45395),
            .in2(N__41781),
            .in3(N__41739),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_16_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_16_13_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_16_13_7  (
            .in0(N__45394),
            .in1(N__45680),
            .in2(N__44829),
            .in3(N__44781),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40320),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_14_1 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_14_1  (
            .in0(N__45980),
            .in1(N__40260),
            .in2(N__41484),
            .in3(N__45406),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_14_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_14_2  (
            .in0(N__45407),
            .in1(N__45981),
            .in2(N__41442),
            .in3(N__40224),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_14_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_14_3  (
            .in0(N__41708),
            .in1(N__45405),
            .in2(N__46012),
            .in3(N__41661),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_14_5 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_16_14_5  (
            .in0(N__45982),
            .in1(N__45404),
            .in2(N__43563),
            .in3(N__43603),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_16_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_16_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_16_14_6  (
            .in0(N__40433),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44576),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_14_7 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_14_7  (
            .in0(N__45976),
            .in1(N__40419),
            .in2(N__41397),
            .in3(N__45408),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_16_15_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_16_15_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_16_15_3  (
            .in0(N__49874),
            .in1(N__42735),
            .in2(N__42204),
            .in3(N__49700),
            .lcout(elapsed_time_ns_1_RNISAHF91_0_13),
            .ltout(elapsed_time_ns_1_RNISAHF91_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_16_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_16_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_16_15_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_16_15_4  (
            .in0(N__40831),
            .in1(N__49574),
            .in2(N__40380),
            .in3(N__46766),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49187),
            .ce(N__48819),
            .sr(N__48419));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_16_15_6 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_16_15_6  (
            .in0(N__42128),
            .in1(N__40365),
            .in2(N__40858),
            .in3(N__46767),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49187),
            .ce(N__48819),
            .sr(N__48419));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_16_0 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_16_16_0  (
            .in0(N__40506),
            .in1(N__43155),
            .in2(N__49876),
            .in3(N__49696),
            .lcout(elapsed_time_ns_1_RNI1HIF91_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_16_1 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_16_16_1  (
            .in0(N__42870),
            .in1(N__40494),
            .in2(N__49711),
            .in3(N__49845),
            .lcout(elapsed_time_ns_1_RNISBIF91_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_16_2 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_16_2  (
            .in0(N__42579),
            .in1(N__49839),
            .in2(N__43227),
            .in3(N__49691),
            .lcout(elapsed_time_ns_1_RNIUDIF91_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_16_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_16_16_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_16_16_3  (
            .in0(N__49690),
            .in1(N__42230),
            .in2(N__49875),
            .in3(N__42759),
            .lcout(elapsed_time_ns_1_RNIR9HF91_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_16_4 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_16_16_4  (
            .in0(N__49840),
            .in1(N__40512),
            .in2(N__43203),
            .in3(N__49692),
            .lcout(elapsed_time_ns_1_RNIVEIF91_0_25),
            .ltout(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_16_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_16_16_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_16_16_5  (
            .in0(N__40481),
            .in1(N__40505),
            .in2(N__40497),
            .in3(N__40469),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_16_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_16_16_6  (
            .in0(N__40493),
            .in1(N__42345),
            .in2(N__40485),
            .in3(N__42567),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_16_7 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_16_16_7  (
            .in0(N__40482),
            .in1(N__49841),
            .in2(N__49710),
            .in3(N__43131),
            .lcout(elapsed_time_ns_1_RNI2IIF91_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_16_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_16_17_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_16_17_0  (
            .in0(N__42105),
            .in1(N__46860),
            .in2(_gnd_net_),
            .in3(N__42158),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_16_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_16_17_1 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_16_17_1  (
            .in0(N__40617),
            .in1(N__49961),
            .in2(N__40635),
            .in3(N__40539),
            .lcout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ),
            .ltout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_17_2 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_16_17_2  (
            .in0(N__40470),
            .in1(N__49701),
            .in2(N__40473),
            .in3(N__43176),
            .lcout(elapsed_time_ns_1_RNI0GIF91_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_17_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_17_3  (
            .in0(N__40458),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47826),
            .lcout(elapsed_time_ns_1_RNIA965M1_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_17_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_17_4  (
            .in0(N__47827),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40452),
            .lcout(elapsed_time_ns_1_RNI9865M1_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_17_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_17_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__42456),
            .in2(_gnd_net_),
            .in3(N__47828),
            .lcout(elapsed_time_ns_1_RNI8765M1_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_17_6 .LUT_INIT=16'b0000110100001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_17_6  (
            .in0(N__40563),
            .in1(N__40545),
            .in2(N__49967),
            .in3(N__42678),
            .lcout(\delay_measurement_inst.delay_tr9 ),
            .ltout(\delay_measurement_inst.delay_tr9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_15_LC_16_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_15_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_15_LC_16_17_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_15_LC_16_17_7  (
            .in0(N__48585),
            .in1(N__40587),
            .in2(N__40548),
            .in3(N__40538),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_21_LC_16_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_21_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_21_LC_16_18_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBSKT4_21_LC_16_18_0  (
            .in0(N__42889),
            .in1(N__42868),
            .in2(_gnd_net_),
            .in3(N__40604),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_17_LC_16_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_17_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_17_LC_16_18_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_17_LC_16_18_1  (
            .in0(N__42714),
            .in1(N__42974),
            .in2(N__42708),
            .in3(N__40596),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_390 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_390_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_17_LC_16_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_17_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_17_LC_16_18_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_17_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40530),
            .in3(N__40631),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_391_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_18_3 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_18_3  (
            .in0(N__48586),
            .in1(N__49962),
            .in2(N__40527),
            .in3(N__40616),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_18_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40524),
            .in3(N__40518),
            .lcout(elapsed_time_ns_1_RNI6565M1_0_14),
            .ltout(elapsed_time_ns_1_RNI6565M1_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_18_5 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_18_5  (
            .in0(N__43068),
            .in1(N__49818),
            .in2(N__40521),
            .in3(N__47615),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_21_LC_16_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_21_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_21_LC_16_18_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_21_LC_16_18_6  (
            .in0(N__42890),
            .in1(N__40605),
            .in2(N__40586),
            .in3(N__42869),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_382 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_382_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_16_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_16_18_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_16_18_7  (
            .in0(N__42696),
            .in1(_gnd_net_),
            .in2(N__40620),
            .in3(N__42442),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_24_LC_16_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_24_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_24_LC_16_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_24_LC_16_19_0  (
            .in0(N__40884),
            .in1(N__43220),
            .in2(N__43199),
            .in3(N__40569),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_356 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_19_2 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_16_19_2  (
            .in0(N__43062),
            .in1(N__46344),
            .in2(N__42829),
            .in3(N__40559),
            .lcout(\delay_measurement_inst.N_363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4DNE1_16_LC_16_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4DNE1_16_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4DNE1_16_LC_16_19_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4DNE1_16_LC_16_19_3  (
            .in0(N__46345),
            .in1(N__47735),
            .in2(N__43007),
            .in3(N__42941),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_19_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_19_4  (
            .in0(N__42728),
            .in1(N__42773),
            .in2(N__42755),
            .in3(N__42791),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_351 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_351_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_15_LC_16_19_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_15_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_15_LC_16_19_5 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_15_LC_16_19_5  (
            .in0(N__43024),
            .in1(_gnd_net_),
            .in2(N__40590),
            .in3(N__42672),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIK0B1_23_LC_16_20_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIK0B1_23_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIK0B1_23_LC_16_20_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIK0B1_23_LC_16_20_3  (
            .in0(N__43088),
            .in1(N__43109),
            .in2(_gnd_net_),
            .in3(N__43241),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_20_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_16_20_5  (
            .in0(N__42940),
            .in1(N__42967),
            .in2(N__43006),
            .in3(N__47728),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_21_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40923),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH8AP1_20_LC_16_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH8AP1_20_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH8AP1_20_LC_16_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH8AP1_20_LC_16_21_5  (
            .in0(N__43124),
            .in1(N__43169),
            .in2(N__43151),
            .in3(N__42908),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_22_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_16_22_1  (
            .in0(N__49576),
            .in1(N__42234),
            .in2(N__40872),
            .in3(N__46822),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49141),
            .ce(N__48820),
            .sr(N__48475));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_16_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_16_22_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_16_22_3  (
            .in0(N__49575),
            .in1(N__46484),
            .in2(_gnd_net_),
            .in3(N__46821),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49141),
            .ce(N__48820),
            .sr(N__48475));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_16_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_16_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_16_22_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_16_22_6  (
            .in0(N__46820),
            .in1(N__47783),
            .in2(_gnd_net_),
            .in3(N__49577),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49141),
            .ce(N__48820),
            .sr(N__48475));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_23_1 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_16_23_1  (
            .in0(N__49578),
            .in1(N__42561),
            .in2(_gnd_net_),
            .in3(N__46819),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49136),
            .ce(N__48801),
            .sr(N__48483));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_5_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_5_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_17_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40733),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49244),
            .ce(N__44136),
            .sr(N__48391));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44898),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_6_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_17_6_1  (
            .in0(N__45424),
            .in1(N__46006),
            .in2(N__40707),
            .in3(N__41252),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40651),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_6_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_17_6_3  (
            .in0(N__45427),
            .in1(N__46004),
            .in2(N__46277),
            .in3(N__46236),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_17_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46269),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_17_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44998),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_6_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_17_6_6  (
            .in0(N__46007),
            .in1(N__45425),
            .in2(N__41102),
            .in3(N__41203),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_6_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_17_6_7  (
            .in0(N__45426),
            .in1(N__46005),
            .in2(N__43700),
            .in3(N__43647),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_7_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(N__43512),
            .in2(N__41056),
            .in3(N__41049),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_7_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_7_1  (
            .in0(_gnd_net_),
            .in1(N__41028),
            .in2(_gnd_net_),
            .in3(N__40998),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_7_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_7_2  (
            .in0(_gnd_net_),
            .in1(N__40995),
            .in2(_gnd_net_),
            .in3(N__40962),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_7_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(N__40959),
            .in2(_gnd_net_),
            .in3(N__40926),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_7_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_7_4  (
            .in0(_gnd_net_),
            .in1(N__41265),
            .in2(_gnd_net_),
            .in3(N__41235),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_7_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_7_5  (
            .in0(_gnd_net_),
            .in1(N__41232),
            .in2(_gnd_net_),
            .in3(N__41220),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_7_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_7_6  (
            .in0(_gnd_net_),
            .in1(N__41217),
            .in2(_gnd_net_),
            .in3(N__41184),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_7_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_7_7  (
            .in0(_gnd_net_),
            .in1(N__41181),
            .in2(_gnd_net_),
            .in3(N__41172),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(N__41169),
            .in2(_gnd_net_),
            .in3(N__41133),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(N__41130),
            .in2(_gnd_net_),
            .in3(N__41124),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(N__41121),
            .in2(_gnd_net_),
            .in3(N__41109),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_8_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43521),
            .in3(N__41106),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(N__41343),
            .in2(_gnd_net_),
            .in3(N__41337),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(N__43344),
            .in2(_gnd_net_),
            .in3(N__41334),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__41331),
            .in2(_gnd_net_),
            .in3(N__41319),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(N__41316),
            .in2(_gnd_net_),
            .in3(N__41307),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__41304),
            .in2(_gnd_net_),
            .in3(N__41295),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__41292),
            .in2(_gnd_net_),
            .in3(N__41283),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__41280),
            .in2(_gnd_net_),
            .in3(N__41271),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__46200),
            .in2(_gnd_net_),
            .in3(N__41268),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__41559),
            .in2(_gnd_net_),
            .in3(N__41538),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(N__41535),
            .in2(_gnd_net_),
            .in3(N__41526),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(N__41523),
            .in2(_gnd_net_),
            .in3(N__41514),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_9_7  (
            .in0(_gnd_net_),
            .in1(N__41511),
            .in2(_gnd_net_),
            .in3(N__41496),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__41493),
            .in2(_gnd_net_),
            .in3(N__41454),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__41451),
            .in2(_gnd_net_),
            .in3(N__41409),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__41406),
            .in2(_gnd_net_),
            .in3(N__41370),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__41367),
            .in2(_gnd_net_),
            .in3(N__41346),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__41796),
            .in2(_gnd_net_),
            .in3(N__41787),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41784),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_10_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_17_10_6  (
            .in0(N__45266),
            .in1(N__45942),
            .in2(N__41780),
            .in3(N__41734),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_17_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_17_10_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_17_10_7  (
            .in0(N__45941),
            .in1(N__45267),
            .in2(N__41709),
            .in3(N__41656),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_17_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_17_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__41637),
            .in2(N__41612),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_17_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_17_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__44093),
            .in2(N__44070),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_17_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_17_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__45888),
            .in2(N__41595),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_17_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_17_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__41586),
            .in2(N__45993),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_17_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_17_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__45892),
            .in2(N__41574),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_17_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_17_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__41847),
            .in2(N__45994),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_17_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_17_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__45896),
            .in2(N__43359),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_17_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_17_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__41838),
            .in2(N__45995),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_17_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_17_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__45751),
            .in2(N__43281),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_17_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_17_12_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__41829),
            .in2(N__45907),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_17_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_17_12_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__45755),
            .in2(N__44757),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_17_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_17_12_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__41817),
            .in2(N__45908),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_17_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_17_12_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__45759),
            .in2(N__41808),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_17_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_17_12_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(N__43440),
            .in2(N__45909),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_17_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_17_12_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__45763),
            .in2(N__46029),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_17_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_17_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__43713),
            .in2(N__45910),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_17_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_17_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__45911),
            .in2(N__43536),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_17_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_17_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__46122),
            .in2(N__45996),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_17_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_17_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__45915),
            .in2(N__44178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_17_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_17_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__44610),
            .in2(N__45997),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_17_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_17_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(N__45919),
            .in2(N__45072),
            .in3(N__41874),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_17_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_17_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__41871),
            .in2(N__45998),
            .in3(N__41850),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_17_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_17_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(N__45923),
            .in2(N__42078),
            .in3(N__42051),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_17_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_17_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(N__44940),
            .in2(N__45999),
            .in3(N__42036),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_17_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_17_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__45927),
            .in2(N__42033),
            .in3(N__42009),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_17_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_17_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__42006),
            .in2(N__46000),
            .in3(N__41988),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_17_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_17_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__45931),
            .in2(N__41985),
            .in3(N__41961),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_17_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_17_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(N__41958),
            .in2(N__46001),
            .in3(N__41934),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_17_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_17_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__45935),
            .in2(N__41931),
            .in3(N__41904),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_17_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_17_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__44841),
            .in2(N__46002),
            .in3(N__41889),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_17_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_17_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(N__45939),
            .in2(N__43869),
            .in3(N__42288),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_17_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_17_14_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_17_14_7  (
            .in0(N__45940),
            .in1(N__45403),
            .in2(_gnd_net_),
            .in3(N__42285),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_17_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_17_15_0 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_17_15_0  (
            .in0(N__49861),
            .in1(N__49686),
            .in2(N__42253),
            .in3(N__42795),
            .lcout(elapsed_time_ns_1_RNIP7HF91_0_10),
            .ltout(elapsed_time_ns_1_RNIP7HF91_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_17_15_1  (
            .in0(N__42225),
            .in1(N__42199),
            .in2(N__42183),
            .in3(N__42321),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_15_2 .LUT_INIT=16'b0011001111110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(N__42169),
            .in2(N__42132),
            .in3(N__42127),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_15_3 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_17_15_3  (
            .in0(N__42388),
            .in1(N__46867),
            .in2(N__42087),
            .in3(N__46727),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_17_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_17_15_4 .LUT_INIT=16'b1111110111101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_17_15_4  (
            .in0(N__49863),
            .in1(N__47842),
            .in2(N__42660),
            .in3(N__46427),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_17_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_17_15_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42084),
            .in3(N__47668),
            .lcout(elapsed_time_ns_1_RNIK8NQL1_0_3),
            .ltout(elapsed_time_ns_1_RNIK8NQL1_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_17_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_17_15_6 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42081),
            .in3(N__46399),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_17_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_17_15_7 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_17_15_7  (
            .in0(N__46400),
            .in1(N__49862),
            .in2(N__49709),
            .in3(N__50013),
            .lcout(elapsed_time_ns_1_RNIAE2591_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_16_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_17_16_0  (
            .in0(N__49679),
            .in1(N__49814),
            .in2(N__42363),
            .in3(N__42894),
            .lcout(elapsed_time_ns_1_RNIRAIF91_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_17_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_17_16_1 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_17_16_1  (
            .in0(N__42449),
            .in1(N__48584),
            .in2(N__42423),
            .in3(N__49951),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_16_2 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_17_16_2  (
            .in0(N__46874),
            .in1(N__43038),
            .in2(N__42414),
            .in3(N__49816),
            .lcout(elapsed_time_ns_1_RNIUCHF91_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_17_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_17_16_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__47841),
            .in2(_gnd_net_),
            .in3(N__47715),
            .lcout(elapsed_time_ns_1_RNIBA65M1_0_19),
            .ltout(elapsed_time_ns_1_RNIBA65M1_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_17_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_17_16_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_17_16_4  (
            .in0(N__42554),
            .in1(N__42515),
            .in2(N__42411),
            .in3(N__46472),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_17_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_17_16_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_17_16_5  (
            .in0(N__49813),
            .in1(N__42372),
            .in2(N__42918),
            .in3(N__49678),
            .lcout(elapsed_time_ns_1_RNIQ9IF91_0_20),
            .ltout(elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_16_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_17_16_6  (
            .in0(N__42599),
            .in1(N__42467),
            .in2(N__42366),
            .in3(N__42356),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_16_7 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_17_16_7  (
            .in0(N__49815),
            .in1(N__42777),
            .in2(N__42335),
            .in3(N__49680),
            .lcout(elapsed_time_ns_1_RNIQ8HF91_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_17_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_17_17_0  (
            .in0(N__49682),
            .in1(N__49820),
            .in2(N__42603),
            .in3(N__43110),
            .lcout(elapsed_time_ns_1_RNI3JIF91_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_17_1 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_17_17_1  (
            .in0(N__49819),
            .in1(N__42588),
            .in2(N__43248),
            .in3(N__49681),
            .lcout(elapsed_time_ns_1_RNITCIF91_0_23),
            .ltout(elapsed_time_ns_1_RNITCIF91_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_17_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42582),
            .in3(N__42578),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_17_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_17_17_3 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_17_17_3  (
            .in0(N__50416),
            .in1(N__42639),
            .in2(N__49864),
            .in3(N__49684),
            .lcout(elapsed_time_ns_1_RNICG2591_0_4),
            .ltout(elapsed_time_ns_1_RNICG2591_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_17_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_17_17_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_17_17_4  (
            .in0(N__47766),
            .in1(N__42555),
            .in2(N__42528),
            .in3(N__46536),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_17_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_17_17_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_17_17_5  (
            .in0(N__42516),
            .in1(N__42485),
            .in2(N__42474),
            .in3(N__46473),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_17_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_17_17_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_17_17_6  (
            .in0(N__49683),
            .in1(N__49821),
            .in2(N__42471),
            .in3(N__43089),
            .lcout(elapsed_time_ns_1_RNIRBJF91_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_17_7 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_17_17_7  (
            .in0(N__46537),
            .in1(N__42621),
            .in2(N__49865),
            .in3(N__49685),
            .lcout(elapsed_time_ns_1_RNIDH2591_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_17_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_17_18_0 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_17_18_0  (
            .in0(N__43008),
            .in1(N__46480),
            .in2(N__49886),
            .in3(N__47626),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_17_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_17_18_2 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_17_18_2  (
            .in0(N__42653),
            .in1(N__50009),
            .in2(N__42830),
            .in3(N__43066),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_17_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_17_18_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__42617),
            .in2(_gnd_net_),
            .in3(N__42635),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_344 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_18_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_17_18_4  (
            .in0(N__42652),
            .in1(N__50008),
            .in2(N__42699),
            .in3(N__50054),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_347 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMF21_6_LC_17_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMF21_6_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMF21_6_LC_17_18_5 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQMF21_6_LC_17_18_5  (
            .in0(N__42825),
            .in1(N__46346),
            .in2(N__42690),
            .in3(N__42671),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID68O3_15_LC_17_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID68O3_15_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID68O3_15_LC_17_18_6 .LUT_INIT=16'b1110111011101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID68O3_15_LC_17_18_6  (
            .in0(N__43037),
            .in1(N__43067),
            .in2(N__42687),
            .in3(N__42684),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_18_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(N__47897),
            .in2(_gnd_net_),
            .in3(N__45032),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_348 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__46594),
            .in2(N__50081),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49165),
            .ce(N__49985),
            .sr(N__48446));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__46570),
            .in2(N__50036),
            .in3(N__42624),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49165),
            .ce(N__49985),
            .sr(N__48446));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(N__47077),
            .in2(N__46599),
            .in3(N__42606),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49165),
            .ce(N__49985),
            .sr(N__48446));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__47053),
            .in2(N__46575),
            .in3(N__42843),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49165),
            .ce(N__49985),
            .sr(N__48446));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__47029),
            .in2(N__47082),
            .in3(N__42840),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49165),
            .ce(N__49985),
            .sr(N__48446));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__47005),
            .in2(N__47058),
            .in3(N__42837),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49165),
            .ce(N__49985),
            .sr(N__48446));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__46981),
            .in2(N__47034),
            .in3(N__42798),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49165),
            .ce(N__49985),
            .sr(N__48446));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(N__46957),
            .in2(N__47010),
            .in3(N__42780),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49165),
            .ce(N__49985),
            .sr(N__48446));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__46933),
            .in2(N__46986),
            .in3(N__42762),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49157),
            .ce(N__49986),
            .sr(N__48456));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__46909),
            .in2(N__46962),
            .in3(N__42738),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49157),
            .ce(N__49986),
            .sr(N__48456));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__47293),
            .in2(N__46938),
            .in3(N__42717),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49157),
            .ce(N__49986),
            .sr(N__48456));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__47269),
            .in2(N__46914),
            .in3(N__43041),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49157),
            .ce(N__49986),
            .sr(N__48456));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__47245),
            .in2(N__47298),
            .in3(N__43011),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49157),
            .ce(N__49986),
            .sr(N__48456));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(N__47221),
            .in2(N__47274),
            .in3(N__42981),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49157),
            .ce(N__49986),
            .sr(N__48456));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__47197),
            .in2(N__47250),
            .in3(N__42951),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49157),
            .ce(N__49986),
            .sr(N__48456));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(N__47173),
            .in2(N__47226),
            .in3(N__42924),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49157),
            .ce(N__49986),
            .sr(N__48456));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(N__47149),
            .in2(N__47202),
            .in3(N__42921),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49152),
            .ce(N__49987),
            .sr(N__48463));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(N__47125),
            .in2(N__47178),
            .in3(N__42897),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49152),
            .ce(N__49987),
            .sr(N__48463));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__47101),
            .in2(N__47154),
            .in3(N__42873),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49152),
            .ce(N__49987),
            .sr(N__48463));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(N__47476),
            .in2(N__47130),
            .in3(N__42846),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49152),
            .ce(N__49987),
            .sr(N__48463));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(N__47452),
            .in2(N__47106),
            .in3(N__43230),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49152),
            .ce(N__49987),
            .sr(N__48463));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(N__47428),
            .in2(N__47481),
            .in3(N__43206),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49152),
            .ce(N__49987),
            .sr(N__48463));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(N__47404),
            .in2(N__47457),
            .in3(N__43179),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49152),
            .ce(N__49987),
            .sr(N__48463));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(N__47380),
            .in2(N__47433),
            .in3(N__43158),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49152),
            .ce(N__49987),
            .sr(N__48463));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(N__47356),
            .in2(N__47409),
            .in3(N__43134),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_17_22_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49147),
            .ce(N__49989),
            .sr(N__48469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_22_1  (
            .in0(_gnd_net_),
            .in1(N__47332),
            .in2(N__47385),
            .in3(N__43113),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49147),
            .ce(N__49989),
            .sr(N__48469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_22_2  (
            .in0(_gnd_net_),
            .in1(N__47312),
            .in2(N__47361),
            .in3(N__43092),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49147),
            .ce(N__49989),
            .sr(N__48469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(N__47957),
            .in2(N__47337),
            .in3(N__43071),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49147),
            .ce(N__49989),
            .sr(N__48469));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_22_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43611),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49147),
            .ce(N__49989),
            .sr(N__48469));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_7_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_18_7_0  (
            .in0(N__46009),
            .in1(N__45431),
            .in2(N__43608),
            .in3(N__43552),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_18_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43693),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_7_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_7_2  (
            .in0(_gnd_net_),
            .in1(N__43914),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_7_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_18_7_4  (
            .in0(N__46008),
            .in1(N__45430),
            .in2(N__43502),
            .in3(N__43457),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_18_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_18_7_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_18_7_5  (
            .in0(N__45428),
            .in1(N__46010),
            .in2(N__43421),
            .in3(N__43378),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46105),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_18_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_18_7_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_18_7_7  (
            .in0(N__45429),
            .in1(N__46011),
            .in2(N__43338),
            .in3(N__43314),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_8_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_8_0  (
            .in0(N__45413),
            .in1(N__43931),
            .in2(N__44103),
            .in3(N__43916),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_8_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44163),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49236),
            .ce(N__44135),
            .sr(N__48392));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_8_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_8_3  (
            .in0(N__43917),
            .in1(N__45414),
            .in2(N__43932),
            .in3(N__44102),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_8_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_8_4  (
            .in0(N__44054),
            .in1(N__43927),
            .in2(_gnd_net_),
            .in3(N__43915),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_8_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(N__45415),
            .in2(_gnd_net_),
            .in3(N__43816),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_8_6 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_8_6  (
            .in0(N__45416),
            .in1(N__43818),
            .in2(N__43854),
            .in3(N__45992),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_8_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_8_7  (
            .in0(N__43850),
            .in1(N__45417),
            .in2(N__46014),
            .in3(N__43817),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_18_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_18_9_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_18_9_0  (
            .in0(N__45954),
            .in1(N__45434),
            .in2(N__43782),
            .in3(N__43732),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_18_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_18_9_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_18_9_1  (
            .in0(N__45433),
            .in1(N__45953),
            .in2(N__43701),
            .in3(N__43646),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_9_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_9_2  (
            .in0(N__45948),
            .in1(N__45436),
            .in2(N__45002),
            .in3(N__44957),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_18_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_18_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_18_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_18_9_3  (
            .in0(_gnd_net_),
            .in1(N__44917),
            .in2(_gnd_net_),
            .in3(N__44589),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_9_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_18_9_4  (
            .in0(N__44899),
            .in1(N__45437),
            .in2(N__46003),
            .in3(N__44857),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_9_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_18_9_5  (
            .in0(N__45432),
            .in1(N__45952),
            .in2(N__44825),
            .in3(N__44774),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_18_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_18_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_18_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_18_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44745),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_9_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_18_9_7  (
            .in0(N__45435),
            .in1(N__45955),
            .in2(N__44675),
            .in3(N__44627),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_18_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_18_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_18_10_0  (
            .in0(N__44588),
            .in1(N__44269),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_18_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_18_10_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_18_10_1  (
            .in0(N__45947),
            .in1(N__45439),
            .in2(N__44243),
            .in3(N__44216),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_18_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_18_10_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_18_10_2  (
            .in0(N__45442),
            .in1(N__45943),
            .in2(N__46281),
            .in3(N__46232),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45101),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_18_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_18_10_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_18_10_5  (
            .in0(N__45946),
            .in1(N__45440),
            .in2(N__46194),
            .in3(N__46139),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_10_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_18_10_6  (
            .in0(N__45438),
            .in1(N__45945),
            .in2(N__46113),
            .in3(N__46052),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_10_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_18_10_7  (
            .in0(N__45944),
            .in1(N__45441),
            .in2(N__45126),
            .in3(N__45102),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_18_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_18_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_18_13_5 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_18_13_5  (
            .in0(N__46428),
            .in1(N__49383),
            .in2(N__46386),
            .in3(N__50384),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49210),
            .ce(N__48821),
            .sr(N__48402));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_18_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_18_15_0 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_18_15_0  (
            .in0(N__49893),
            .in1(N__47527),
            .in2(N__45042),
            .in3(N__49705),
            .lcout(elapsed_time_ns_1_RNIFJ2591_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_18_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_18_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_18_15_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_18_15_3  (
            .in0(N__50348),
            .in1(N__49538),
            .in2(_gnd_net_),
            .in3(N__47885),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49199),
            .ce(N__50284),
            .sr(N__48407));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_18_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_18_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_18_15_4 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_18_15_4  (
            .in0(N__49367),
            .in1(N__50349),
            .in2(N__49579),
            .in3(N__46547),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49199),
            .ce(N__50284),
            .sr(N__48407));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_18_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_18_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_18_15_5 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_18_15_5  (
            .in0(N__46382),
            .in1(N__49368),
            .in2(N__50383),
            .in3(N__46423),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49199),
            .ce(N__50284),
            .sr(N__48407));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_18_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_18_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_18_15_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_18_15_6  (
            .in0(N__49537),
            .in1(N__46485),
            .in2(_gnd_net_),
            .in3(N__46818),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49199),
            .ce(N__50284),
            .sr(N__48407));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_18_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_18_16_0 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_18_16_0  (
            .in0(N__46368),
            .in1(N__46422),
            .in2(N__46299),
            .in3(N__46401),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_18_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_18_16_1 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_18_16_1  (
            .in0(N__49464),
            .in1(N__46294),
            .in2(N__46808),
            .in3(N__46367),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_18_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_18_16_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_18_16_2  (
            .in0(N__46366),
            .in1(N__46772),
            .in2(N__46298),
            .in3(N__46356),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_18_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_18_16_3 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_18_16_3  (
            .in0(N__47662),
            .in1(N__46630),
            .in2(N__49905),
            .in3(N__46350),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_18_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_18_16_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46326),
            .in3(N__47846),
            .lcout(elapsed_time_ns_1_RNINBNQL1_0_6),
            .ltout(elapsed_time_ns_1_RNINBNQL1_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_18_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_18_16_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_18_16_5  (
            .in0(N__47881),
            .in1(N__47520),
            .in2(N__46323),
            .in3(N__46310),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_18_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_18_16_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__46868),
            .in2(N__46827),
            .in3(N__46768),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_18_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_18_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_18_16_7 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_18_16_7  (
            .in0(N__49465),
            .in1(N__46631),
            .in2(N__46671),
            .in3(N__50385),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49194),
            .ce(N__50280),
            .sr(N__48414));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_0 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_18_17_0  (
            .in0(N__49364),
            .in1(N__50394),
            .in2(N__49607),
            .in3(N__50420),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49188),
            .ce(N__48811),
            .sr(N__48420));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_18_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_18_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_18_17_3 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_18_17_3  (
            .in0(N__50447),
            .in1(N__49366),
            .in2(N__50400),
            .in3(N__49606),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49188),
            .ce(N__48811),
            .sr(N__48420));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_18_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_18_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_18_17_6 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_18_17_6  (
            .in0(N__49365),
            .in1(N__50395),
            .in2(N__49608),
            .in3(N__46632),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49188),
            .ce(N__48811),
            .sr(N__48420));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_18_18_0  (
            .in0(N__48083),
            .in1(N__50074),
            .in2(_gnd_net_),
            .in3(N__46605),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__49181),
            .ce(N__47934),
            .sr(N__48429));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_18_18_1  (
            .in0(N__48061),
            .in1(N__50029),
            .in2(_gnd_net_),
            .in3(N__46602),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__49181),
            .ce(N__47934),
            .sr(N__48429));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_18_18_2  (
            .in0(N__48084),
            .in1(N__46595),
            .in2(_gnd_net_),
            .in3(N__46578),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__49181),
            .ce(N__47934),
            .sr(N__48429));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_18_18_3  (
            .in0(N__48062),
            .in1(N__46571),
            .in2(_gnd_net_),
            .in3(N__46554),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__49181),
            .ce(N__47934),
            .sr(N__48429));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_18_18_4  (
            .in0(N__48085),
            .in1(N__47078),
            .in2(_gnd_net_),
            .in3(N__47061),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__49181),
            .ce(N__47934),
            .sr(N__48429));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_18_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_18_18_5  (
            .in0(N__48063),
            .in1(N__47054),
            .in2(_gnd_net_),
            .in3(N__47037),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__49181),
            .ce(N__47934),
            .sr(N__48429));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_18_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_18_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_18_18_6  (
            .in0(N__48086),
            .in1(N__47030),
            .in2(_gnd_net_),
            .in3(N__47013),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__49181),
            .ce(N__47934),
            .sr(N__48429));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_18_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_18_18_7  (
            .in0(N__48064),
            .in1(N__47006),
            .in2(_gnd_net_),
            .in3(N__46989),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__49181),
            .ce(N__47934),
            .sr(N__48429));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_18_19_0  (
            .in0(N__48068),
            .in1(N__46982),
            .in2(_gnd_net_),
            .in3(N__46965),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__49173),
            .ce(N__47945),
            .sr(N__48435));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_18_19_1  (
            .in0(N__48076),
            .in1(N__46958),
            .in2(_gnd_net_),
            .in3(N__46941),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__49173),
            .ce(N__47945),
            .sr(N__48435));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_18_19_2  (
            .in0(N__48065),
            .in1(N__46934),
            .in2(_gnd_net_),
            .in3(N__46917),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__49173),
            .ce(N__47945),
            .sr(N__48435));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_18_19_3  (
            .in0(N__48073),
            .in1(N__46910),
            .in2(_gnd_net_),
            .in3(N__46893),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__49173),
            .ce(N__47945),
            .sr(N__48435));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_18_19_4  (
            .in0(N__48066),
            .in1(N__47294),
            .in2(_gnd_net_),
            .in3(N__47277),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__49173),
            .ce(N__47945),
            .sr(N__48435));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_18_19_5  (
            .in0(N__48074),
            .in1(N__47270),
            .in2(_gnd_net_),
            .in3(N__47253),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__49173),
            .ce(N__47945),
            .sr(N__48435));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_18_19_6  (
            .in0(N__48067),
            .in1(N__47246),
            .in2(_gnd_net_),
            .in3(N__47229),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__49173),
            .ce(N__47945),
            .sr(N__48435));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_18_19_7  (
            .in0(N__48075),
            .in1(N__47222),
            .in2(_gnd_net_),
            .in3(N__47205),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__49173),
            .ce(N__47945),
            .sr(N__48435));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_18_20_0  (
            .in0(N__48087),
            .in1(N__47198),
            .in2(_gnd_net_),
            .in3(N__47181),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__49166),
            .ce(N__47944),
            .sr(N__48447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_18_20_1  (
            .in0(N__48069),
            .in1(N__47174),
            .in2(_gnd_net_),
            .in3(N__47157),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__49166),
            .ce(N__47944),
            .sr(N__48447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_18_20_2  (
            .in0(N__48088),
            .in1(N__47150),
            .in2(_gnd_net_),
            .in3(N__47133),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__49166),
            .ce(N__47944),
            .sr(N__48447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_18_20_3  (
            .in0(N__48070),
            .in1(N__47126),
            .in2(_gnd_net_),
            .in3(N__47109),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__49166),
            .ce(N__47944),
            .sr(N__48447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_20_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_18_20_4  (
            .in0(N__48089),
            .in1(N__47102),
            .in2(_gnd_net_),
            .in3(N__47085),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__49166),
            .ce(N__47944),
            .sr(N__48447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_20_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_20_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_18_20_5  (
            .in0(N__48071),
            .in1(N__47477),
            .in2(_gnd_net_),
            .in3(N__47460),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__49166),
            .ce(N__47944),
            .sr(N__48447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_20_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_18_20_6  (
            .in0(N__48090),
            .in1(N__47453),
            .in2(_gnd_net_),
            .in3(N__47436),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__49166),
            .ce(N__47944),
            .sr(N__48447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_20_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_20_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_18_20_7  (
            .in0(N__48072),
            .in1(N__47429),
            .in2(_gnd_net_),
            .in3(N__47412),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__49166),
            .ce(N__47944),
            .sr(N__48447));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_18_21_0  (
            .in0(N__48077),
            .in1(N__47405),
            .in2(_gnd_net_),
            .in3(N__47388),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__49158),
            .ce(N__47946),
            .sr(N__48457));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_18_21_1  (
            .in0(N__48081),
            .in1(N__47381),
            .in2(_gnd_net_),
            .in3(N__47364),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__49158),
            .ce(N__47946),
            .sr(N__48457));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_18_21_2  (
            .in0(N__48078),
            .in1(N__47357),
            .in2(_gnd_net_),
            .in3(N__47340),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__49158),
            .ce(N__47946),
            .sr(N__48457));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_18_21_3  (
            .in0(N__48082),
            .in1(N__47333),
            .in2(_gnd_net_),
            .in3(N__47316),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__49158),
            .ce(N__47946),
            .sr(N__48457));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_18_21_4  (
            .in0(N__48079),
            .in1(N__47313),
            .in2(_gnd_net_),
            .in3(N__47301),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__49158),
            .ce(N__47946),
            .sr(N__48457));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_21_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_21_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_18_21_5  (
            .in0(N__47958),
            .in1(N__48080),
            .in2(_gnd_net_),
            .in3(N__47961),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49158),
            .ce(N__47946),
            .sr(N__48457));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_20_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_20_13_4 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_20_13_4  (
            .in0(N__47871),
            .in1(N__49900),
            .in2(N__47907),
            .in3(N__49716),
            .lcout(elapsed_time_ns_1_RNIGK2591_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_20_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_20_15_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_20_15_0  (
            .in0(_gnd_net_),
            .in1(N__47544),
            .in2(_gnd_net_),
            .in3(N__47847),
            .lcout(elapsed_time_ns_1_RNII6NQL1_0_1),
            .ltout(elapsed_time_ns_1_RNII6NQL1_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_20_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_20_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_20_15_1 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_20_15_1  (
            .in0(N__49451),
            .in1(_gnd_net_),
            .in2(N__47787),
            .in3(N__50359),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_20_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_20_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_20_15_6 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_20_15_6  (
            .in0(N__47782),
            .in1(N__49888),
            .in2(N__47701),
            .in3(N__47742),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_20_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_20_15_7 .LUT_INIT=16'b1111111101001110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_20_15_7  (
            .in0(N__49889),
            .in1(N__49315),
            .in2(N__50058),
            .in3(N__47690),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_20_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_20_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_20_16_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_20_16_0  (
            .in0(N__47537),
            .in1(N__49458),
            .in2(_gnd_net_),
            .in3(N__50391),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49205),
            .ce(N__50286),
            .sr(N__48415));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_20_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_20_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_20_16_3 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_20_16_3  (
            .in0(N__49372),
            .in1(N__49316),
            .in2(N__49281),
            .in3(N__49298),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49205),
            .ce(N__50286),
            .sr(N__48415));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_20_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_20_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_20_16_6 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_20_16_6  (
            .in0(N__50451),
            .in1(N__49374),
            .in2(N__50399),
            .in3(N__49459),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49205),
            .ce(N__50286),
            .sr(N__48415));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_20_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_20_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_20_16_7 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_20_16_7  (
            .in0(N__49373),
            .in1(N__49460),
            .in2(N__50427),
            .in3(N__50390),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49205),
            .ce(N__50286),
            .sr(N__48415));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_20_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50082),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49195),
            .ce(N__49988),
            .sr(N__48430));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_20_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_20_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_20_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_20_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50037),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49195),
            .ce(N__49988),
            .sr(N__48430));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_21_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_21_16_3 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_21_16_3  (
            .in0(N__49963),
            .in1(N__49904),
            .in2(N__49498),
            .in3(N__49715),
            .lcout(elapsed_time_ns_1_RNISCJF91_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_21_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_21_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_21_16_5 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_21_16_5  (
            .in0(N__49381),
            .in1(N__49317),
            .in2(N__49299),
            .in3(N__49280),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49212),
            .ce(N__48822),
            .sr(N__48421));
endmodule // MAIN
