// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 14 2025 21:01:10

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_g,
    T01,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_g;
    output T01;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__50557;
    wire N__50556;
    wire N__50555;
    wire N__50546;
    wire N__50545;
    wire N__50544;
    wire N__50537;
    wire N__50536;
    wire N__50535;
    wire N__50528;
    wire N__50527;
    wire N__50526;
    wire N__50519;
    wire N__50518;
    wire N__50517;
    wire N__50510;
    wire N__50509;
    wire N__50508;
    wire N__50501;
    wire N__50500;
    wire N__50499;
    wire N__50492;
    wire N__50491;
    wire N__50490;
    wire N__50483;
    wire N__50482;
    wire N__50481;
    wire N__50474;
    wire N__50473;
    wire N__50472;
    wire N__50465;
    wire N__50464;
    wire N__50463;
    wire N__50456;
    wire N__50455;
    wire N__50454;
    wire N__50447;
    wire N__50446;
    wire N__50445;
    wire N__50438;
    wire N__50437;
    wire N__50436;
    wire N__50429;
    wire N__50428;
    wire N__50427;
    wire N__50420;
    wire N__50419;
    wire N__50418;
    wire N__50411;
    wire N__50410;
    wire N__50409;
    wire N__50392;
    wire N__50391;
    wire N__50388;
    wire N__50385;
    wire N__50380;
    wire N__50379;
    wire N__50376;
    wire N__50373;
    wire N__50370;
    wire N__50365;
    wire N__50362;
    wire N__50359;
    wire N__50358;
    wire N__50355;
    wire N__50352;
    wire N__50349;
    wire N__50344;
    wire N__50343;
    wire N__50340;
    wire N__50337;
    wire N__50334;
    wire N__50329;
    wire N__50326;
    wire N__50323;
    wire N__50322;
    wire N__50321;
    wire N__50320;
    wire N__50317;
    wire N__50314;
    wire N__50311;
    wire N__50308;
    wire N__50307;
    wire N__50306;
    wire N__50305;
    wire N__50304;
    wire N__50303;
    wire N__50302;
    wire N__50301;
    wire N__50296;
    wire N__50295;
    wire N__50294;
    wire N__50293;
    wire N__50292;
    wire N__50291;
    wire N__50290;
    wire N__50289;
    wire N__50288;
    wire N__50285;
    wire N__50284;
    wire N__50283;
    wire N__50282;
    wire N__50281;
    wire N__50280;
    wire N__50279;
    wire N__50278;
    wire N__50277;
    wire N__50276;
    wire N__50275;
    wire N__50274;
    wire N__50273;
    wire N__50272;
    wire N__50271;
    wire N__50270;
    wire N__50269;
    wire N__50266;
    wire N__50259;
    wire N__50250;
    wire N__50247;
    wire N__50240;
    wire N__50237;
    wire N__50228;
    wire N__50225;
    wire N__50216;
    wire N__50207;
    wire N__50198;
    wire N__50189;
    wire N__50184;
    wire N__50181;
    wire N__50172;
    wire N__50165;
    wire N__50160;
    wire N__50155;
    wire N__50152;
    wire N__50149;
    wire N__50140;
    wire N__50139;
    wire N__50136;
    wire N__50133;
    wire N__50132;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50112;
    wire N__50107;
    wire N__50106;
    wire N__50103;
    wire N__50102;
    wire N__50099;
    wire N__50098;
    wire N__50095;
    wire N__50092;
    wire N__50089;
    wire N__50088;
    wire N__50085;
    wire N__50082;
    wire N__50079;
    wire N__50076;
    wire N__50073;
    wire N__50062;
    wire N__50059;
    wire N__50058;
    wire N__50055;
    wire N__50052;
    wire N__50049;
    wire N__50046;
    wire N__50041;
    wire N__50038;
    wire N__50037;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50025;
    wire N__50022;
    wire N__50019;
    wire N__50018;
    wire N__50017;
    wire N__50016;
    wire N__50011;
    wire N__50006;
    wire N__50003;
    wire N__49998;
    wire N__49993;
    wire N__49990;
    wire N__49989;
    wire N__49986;
    wire N__49983;
    wire N__49978;
    wire N__49977;
    wire N__49976;
    wire N__49975;
    wire N__49974;
    wire N__49973;
    wire N__49972;
    wire N__49971;
    wire N__49970;
    wire N__49969;
    wire N__49968;
    wire N__49967;
    wire N__49966;
    wire N__49965;
    wire N__49964;
    wire N__49963;
    wire N__49962;
    wire N__49961;
    wire N__49960;
    wire N__49959;
    wire N__49958;
    wire N__49957;
    wire N__49956;
    wire N__49955;
    wire N__49954;
    wire N__49953;
    wire N__49952;
    wire N__49951;
    wire N__49950;
    wire N__49949;
    wire N__49948;
    wire N__49947;
    wire N__49946;
    wire N__49945;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49941;
    wire N__49940;
    wire N__49939;
    wire N__49938;
    wire N__49937;
    wire N__49936;
    wire N__49935;
    wire N__49934;
    wire N__49933;
    wire N__49932;
    wire N__49931;
    wire N__49930;
    wire N__49929;
    wire N__49928;
    wire N__49927;
    wire N__49926;
    wire N__49925;
    wire N__49924;
    wire N__49923;
    wire N__49922;
    wire N__49921;
    wire N__49920;
    wire N__49919;
    wire N__49918;
    wire N__49917;
    wire N__49916;
    wire N__49915;
    wire N__49914;
    wire N__49913;
    wire N__49912;
    wire N__49911;
    wire N__49910;
    wire N__49909;
    wire N__49908;
    wire N__49907;
    wire N__49906;
    wire N__49905;
    wire N__49904;
    wire N__49903;
    wire N__49902;
    wire N__49901;
    wire N__49900;
    wire N__49899;
    wire N__49898;
    wire N__49897;
    wire N__49896;
    wire N__49895;
    wire N__49894;
    wire N__49893;
    wire N__49892;
    wire N__49891;
    wire N__49890;
    wire N__49889;
    wire N__49888;
    wire N__49887;
    wire N__49886;
    wire N__49885;
    wire N__49884;
    wire N__49883;
    wire N__49882;
    wire N__49881;
    wire N__49880;
    wire N__49879;
    wire N__49878;
    wire N__49877;
    wire N__49876;
    wire N__49875;
    wire N__49874;
    wire N__49873;
    wire N__49872;
    wire N__49871;
    wire N__49870;
    wire N__49869;
    wire N__49868;
    wire N__49867;
    wire N__49866;
    wire N__49865;
    wire N__49864;
    wire N__49863;
    wire N__49862;
    wire N__49861;
    wire N__49860;
    wire N__49859;
    wire N__49858;
    wire N__49857;
    wire N__49856;
    wire N__49855;
    wire N__49854;
    wire N__49853;
    wire N__49852;
    wire N__49851;
    wire N__49850;
    wire N__49591;
    wire N__49588;
    wire N__49587;
    wire N__49586;
    wire N__49585;
    wire N__49584;
    wire N__49583;
    wire N__49582;
    wire N__49581;
    wire N__49580;
    wire N__49577;
    wire N__49574;
    wire N__49571;
    wire N__49568;
    wire N__49565;
    wire N__49562;
    wire N__49559;
    wire N__49554;
    wire N__49551;
    wire N__49548;
    wire N__49545;
    wire N__49544;
    wire N__49543;
    wire N__49542;
    wire N__49541;
    wire N__49540;
    wire N__49539;
    wire N__49538;
    wire N__49537;
    wire N__49536;
    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49532;
    wire N__49531;
    wire N__49530;
    wire N__49529;
    wire N__49528;
    wire N__49527;
    wire N__49526;
    wire N__49525;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49521;
    wire N__49520;
    wire N__49519;
    wire N__49518;
    wire N__49517;
    wire N__49516;
    wire N__49515;
    wire N__49514;
    wire N__49513;
    wire N__49512;
    wire N__49511;
    wire N__49510;
    wire N__49509;
    wire N__49508;
    wire N__49507;
    wire N__49506;
    wire N__49505;
    wire N__49504;
    wire N__49503;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49499;
    wire N__49498;
    wire N__49497;
    wire N__49496;
    wire N__49495;
    wire N__49494;
    wire N__49493;
    wire N__49492;
    wire N__49491;
    wire N__49490;
    wire N__49489;
    wire N__49488;
    wire N__49487;
    wire N__49486;
    wire N__49485;
    wire N__49484;
    wire N__49483;
    wire N__49482;
    wire N__49481;
    wire N__49480;
    wire N__49479;
    wire N__49478;
    wire N__49475;
    wire N__49474;
    wire N__49473;
    wire N__49472;
    wire N__49471;
    wire N__49470;
    wire N__49469;
    wire N__49468;
    wire N__49467;
    wire N__49466;
    wire N__49465;
    wire N__49464;
    wire N__49463;
    wire N__49462;
    wire N__49461;
    wire N__49460;
    wire N__49459;
    wire N__49458;
    wire N__49457;
    wire N__49456;
    wire N__49453;
    wire N__49452;
    wire N__49451;
    wire N__49450;
    wire N__49449;
    wire N__49448;
    wire N__49445;
    wire N__49444;
    wire N__49443;
    wire N__49442;
    wire N__49441;
    wire N__49440;
    wire N__49439;
    wire N__49438;
    wire N__49437;
    wire N__49436;
    wire N__49435;
    wire N__49434;
    wire N__49433;
    wire N__49432;
    wire N__49431;
    wire N__49430;
    wire N__49427;
    wire N__49426;
    wire N__49425;
    wire N__49424;
    wire N__49423;
    wire N__49422;
    wire N__49421;
    wire N__49420;
    wire N__49417;
    wire N__49416;
    wire N__49415;
    wire N__49414;
    wire N__49413;
    wire N__49412;
    wire N__49411;
    wire N__49410;
    wire N__49409;
    wire N__49408;
    wire N__49407;
    wire N__49406;
    wire N__49405;
    wire N__49138;
    wire N__49135;
    wire N__49132;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49122;
    wire N__49121;
    wire N__49120;
    wire N__49117;
    wire N__49114;
    wire N__49111;
    wire N__49110;
    wire N__49109;
    wire N__49108;
    wire N__49105;
    wire N__49104;
    wire N__49103;
    wire N__49102;
    wire N__49101;
    wire N__49100;
    wire N__49099;
    wire N__49098;
    wire N__49095;
    wire N__49094;
    wire N__49093;
    wire N__49092;
    wire N__49091;
    wire N__49090;
    wire N__49089;
    wire N__49088;
    wire N__49087;
    wire N__49086;
    wire N__49085;
    wire N__49084;
    wire N__49083;
    wire N__49082;
    wire N__49081;
    wire N__49080;
    wire N__49079;
    wire N__49076;
    wire N__49073;
    wire N__49070;
    wire N__49069;
    wire N__49066;
    wire N__49063;
    wire N__49060;
    wire N__49051;
    wire N__49044;
    wire N__49041;
    wire N__49032;
    wire N__49023;
    wire N__49014;
    wire N__49005;
    wire N__48998;
    wire N__48995;
    wire N__48994;
    wire N__48993;
    wire N__48990;
    wire N__48987;
    wire N__48986;
    wire N__48985;
    wire N__48984;
    wire N__48983;
    wire N__48980;
    wire N__48975;
    wire N__48964;
    wire N__48963;
    wire N__48962;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48952;
    wire N__48951;
    wire N__48948;
    wire N__48943;
    wire N__48934;
    wire N__48929;
    wire N__48926;
    wire N__48919;
    wire N__48912;
    wire N__48909;
    wire N__48896;
    wire N__48893;
    wire N__48888;
    wire N__48883;
    wire N__48880;
    wire N__48877;
    wire N__48876;
    wire N__48873;
    wire N__48870;
    wire N__48867;
    wire N__48862;
    wire N__48861;
    wire N__48858;
    wire N__48855;
    wire N__48852;
    wire N__48847;
    wire N__48844;
    wire N__48841;
    wire N__48838;
    wire N__48835;
    wire N__48832;
    wire N__48831;
    wire N__48828;
    wire N__48825;
    wire N__48820;
    wire N__48819;
    wire N__48816;
    wire N__48813;
    wire N__48808;
    wire N__48805;
    wire N__48802;
    wire N__48801;
    wire N__48798;
    wire N__48795;
    wire N__48792;
    wire N__48787;
    wire N__48786;
    wire N__48783;
    wire N__48780;
    wire N__48777;
    wire N__48772;
    wire N__48769;
    wire N__48766;
    wire N__48765;
    wire N__48762;
    wire N__48759;
    wire N__48754;
    wire N__48753;
    wire N__48750;
    wire N__48747;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48735;
    wire N__48734;
    wire N__48731;
    wire N__48728;
    wire N__48725;
    wire N__48722;
    wire N__48715;
    wire N__48712;
    wire N__48711;
    wire N__48710;
    wire N__48707;
    wire N__48706;
    wire N__48703;
    wire N__48700;
    wire N__48697;
    wire N__48694;
    wire N__48691;
    wire N__48686;
    wire N__48679;
    wire N__48676;
    wire N__48673;
    wire N__48670;
    wire N__48669;
    wire N__48666;
    wire N__48665;
    wire N__48662;
    wire N__48659;
    wire N__48656;
    wire N__48651;
    wire N__48648;
    wire N__48643;
    wire N__48640;
    wire N__48637;
    wire N__48634;
    wire N__48631;
    wire N__48628;
    wire N__48625;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48615;
    wire N__48612;
    wire N__48609;
    wire N__48606;
    wire N__48601;
    wire N__48598;
    wire N__48595;
    wire N__48594;
    wire N__48591;
    wire N__48588;
    wire N__48585;
    wire N__48580;
    wire N__48577;
    wire N__48576;
    wire N__48573;
    wire N__48570;
    wire N__48567;
    wire N__48562;
    wire N__48559;
    wire N__48558;
    wire N__48555;
    wire N__48552;
    wire N__48549;
    wire N__48544;
    wire N__48541;
    wire N__48540;
    wire N__48537;
    wire N__48534;
    wire N__48531;
    wire N__48526;
    wire N__48523;
    wire N__48520;
    wire N__48519;
    wire N__48514;
    wire N__48513;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48499;
    wire N__48496;
    wire N__48495;
    wire N__48494;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48478;
    wire N__48475;
    wire N__48474;
    wire N__48471;
    wire N__48468;
    wire N__48467;
    wire N__48464;
    wire N__48461;
    wire N__48458;
    wire N__48455;
    wire N__48452;
    wire N__48445;
    wire N__48442;
    wire N__48439;
    wire N__48436;
    wire N__48435;
    wire N__48432;
    wire N__48429;
    wire N__48426;
    wire N__48423;
    wire N__48418;
    wire N__48415;
    wire N__48414;
    wire N__48411;
    wire N__48408;
    wire N__48405;
    wire N__48400;
    wire N__48397;
    wire N__48396;
    wire N__48393;
    wire N__48390;
    wire N__48387;
    wire N__48382;
    wire N__48379;
    wire N__48378;
    wire N__48375;
    wire N__48372;
    wire N__48369;
    wire N__48364;
    wire N__48361;
    wire N__48360;
    wire N__48357;
    wire N__48354;
    wire N__48351;
    wire N__48346;
    wire N__48343;
    wire N__48342;
    wire N__48339;
    wire N__48336;
    wire N__48333;
    wire N__48328;
    wire N__48325;
    wire N__48324;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48303;
    wire N__48300;
    wire N__48297;
    wire N__48294;
    wire N__48289;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48279;
    wire N__48276;
    wire N__48273;
    wire N__48270;
    wire N__48265;
    wire N__48262;
    wire N__48261;
    wire N__48258;
    wire N__48255;
    wire N__48250;
    wire N__48247;
    wire N__48246;
    wire N__48243;
    wire N__48240;
    wire N__48235;
    wire N__48232;
    wire N__48231;
    wire N__48228;
    wire N__48225;
    wire N__48220;
    wire N__48217;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48205;
    wire N__48202;
    wire N__48201;
    wire N__48200;
    wire N__48197;
    wire N__48194;
    wire N__48191;
    wire N__48184;
    wire N__48181;
    wire N__48178;
    wire N__48175;
    wire N__48172;
    wire N__48171;
    wire N__48170;
    wire N__48167;
    wire N__48166;
    wire N__48163;
    wire N__48160;
    wire N__48157;
    wire N__48154;
    wire N__48151;
    wire N__48142;
    wire N__48141;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48124;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48114;
    wire N__48111;
    wire N__48108;
    wire N__48105;
    wire N__48100;
    wire N__48097;
    wire N__48094;
    wire N__48093;
    wire N__48088;
    wire N__48087;
    wire N__48084;
    wire N__48081;
    wire N__48078;
    wire N__48073;
    wire N__48070;
    wire N__48069;
    wire N__48064;
    wire N__48063;
    wire N__48060;
    wire N__48057;
    wire N__48054;
    wire N__48049;
    wire N__48046;
    wire N__48043;
    wire N__48042;
    wire N__48037;
    wire N__48036;
    wire N__48033;
    wire N__48030;
    wire N__48027;
    wire N__48022;
    wire N__48019;
    wire N__48016;
    wire N__48013;
    wire N__48010;
    wire N__48009;
    wire N__48006;
    wire N__48003;
    wire N__48000;
    wire N__47995;
    wire N__47992;
    wire N__47989;
    wire N__47986;
    wire N__47985;
    wire N__47982;
    wire N__47979;
    wire N__47976;
    wire N__47971;
    wire N__47968;
    wire N__47965;
    wire N__47962;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47952;
    wire N__47947;
    wire N__47944;
    wire N__47941;
    wire N__47940;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47926;
    wire N__47923;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47908;
    wire N__47905;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47895;
    wire N__47890;
    wire N__47887;
    wire N__47886;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47872;
    wire N__47869;
    wire N__47868;
    wire N__47865;
    wire N__47862;
    wire N__47859;
    wire N__47854;
    wire N__47851;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47836;
    wire N__47833;
    wire N__47832;
    wire N__47829;
    wire N__47826;
    wire N__47823;
    wire N__47818;
    wire N__47815;
    wire N__47814;
    wire N__47813;
    wire N__47808;
    wire N__47805;
    wire N__47802;
    wire N__47797;
    wire N__47794;
    wire N__47793;
    wire N__47792;
    wire N__47791;
    wire N__47786;
    wire N__47781;
    wire N__47776;
    wire N__47775;
    wire N__47772;
    wire N__47767;
    wire N__47764;
    wire N__47763;
    wire N__47762;
    wire N__47759;
    wire N__47756;
    wire N__47753;
    wire N__47746;
    wire N__47743;
    wire N__47742;
    wire N__47739;
    wire N__47738;
    wire N__47735;
    wire N__47734;
    wire N__47731;
    wire N__47724;
    wire N__47719;
    wire N__47718;
    wire N__47715;
    wire N__47712;
    wire N__47711;
    wire N__47708;
    wire N__47705;
    wire N__47702;
    wire N__47697;
    wire N__47694;
    wire N__47689;
    wire N__47686;
    wire N__47683;
    wire N__47680;
    wire N__47679;
    wire N__47676;
    wire N__47673;
    wire N__47670;
    wire N__47669;
    wire N__47664;
    wire N__47661;
    wire N__47656;
    wire N__47655;
    wire N__47652;
    wire N__47649;
    wire N__47646;
    wire N__47641;
    wire N__47638;
    wire N__47635;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47623;
    wire N__47622;
    wire N__47619;
    wire N__47616;
    wire N__47613;
    wire N__47608;
    wire N__47605;
    wire N__47602;
    wire N__47601;
    wire N__47598;
    wire N__47595;
    wire N__47592;
    wire N__47587;
    wire N__47584;
    wire N__47583;
    wire N__47580;
    wire N__47577;
    wire N__47574;
    wire N__47569;
    wire N__47566;
    wire N__47565;
    wire N__47562;
    wire N__47559;
    wire N__47556;
    wire N__47551;
    wire N__47548;
    wire N__47545;
    wire N__47544;
    wire N__47541;
    wire N__47538;
    wire N__47535;
    wire N__47530;
    wire N__47527;
    wire N__47526;
    wire N__47523;
    wire N__47520;
    wire N__47517;
    wire N__47512;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47498;
    wire N__47495;
    wire N__47492;
    wire N__47489;
    wire N__47486;
    wire N__47479;
    wire N__47478;
    wire N__47477;
    wire N__47476;
    wire N__47475;
    wire N__47464;
    wire N__47461;
    wire N__47458;
    wire N__47455;
    wire N__47452;
    wire N__47451;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47433;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47421;
    wire N__47418;
    wire N__47415;
    wire N__47410;
    wire N__47407;
    wire N__47406;
    wire N__47403;
    wire N__47400;
    wire N__47395;
    wire N__47392;
    wire N__47389;
    wire N__47386;
    wire N__47383;
    wire N__47382;
    wire N__47381;
    wire N__47378;
    wire N__47373;
    wire N__47368;
    wire N__47365;
    wire N__47364;
    wire N__47361;
    wire N__47358;
    wire N__47355;
    wire N__47352;
    wire N__47351;
    wire N__47348;
    wire N__47345;
    wire N__47342;
    wire N__47335;
    wire N__47332;
    wire N__47329;
    wire N__47326;
    wire N__47323;
    wire N__47322;
    wire N__47319;
    wire N__47316;
    wire N__47311;
    wire N__47308;
    wire N__47305;
    wire N__47302;
    wire N__47299;
    wire N__47296;
    wire N__47293;
    wire N__47292;
    wire N__47291;
    wire N__47288;
    wire N__47285;
    wire N__47282;
    wire N__47275;
    wire N__47272;
    wire N__47269;
    wire N__47266;
    wire N__47265;
    wire N__47264;
    wire N__47261;
    wire N__47258;
    wire N__47255;
    wire N__47248;
    wire N__47245;
    wire N__47242;
    wire N__47239;
    wire N__47236;
    wire N__47233;
    wire N__47230;
    wire N__47227;
    wire N__47226;
    wire N__47225;
    wire N__47222;
    wire N__47217;
    wire N__47212;
    wire N__47209;
    wire N__47208;
    wire N__47207;
    wire N__47204;
    wire N__47199;
    wire N__47194;
    wire N__47193;
    wire N__47190;
    wire N__47189;
    wire N__47186;
    wire N__47183;
    wire N__47180;
    wire N__47173;
    wire N__47172;
    wire N__47171;
    wire N__47168;
    wire N__47163;
    wire N__47160;
    wire N__47157;
    wire N__47152;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47128;
    wire N__47125;
    wire N__47124;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47112;
    wire N__47111;
    wire N__47108;
    wire N__47107;
    wire N__47106;
    wire N__47105;
    wire N__47102;
    wire N__47099;
    wire N__47098;
    wire N__47097;
    wire N__47094;
    wire N__47089;
    wire N__47088;
    wire N__47087;
    wire N__47086;
    wire N__47085;
    wire N__47084;
    wire N__47083;
    wire N__47080;
    wire N__47079;
    wire N__47078;
    wire N__47077;
    wire N__47076;
    wire N__47073;
    wire N__47072;
    wire N__47071;
    wire N__47070;
    wire N__47069;
    wire N__47068;
    wire N__47067;
    wire N__47066;
    wire N__47065;
    wire N__47064;
    wire N__47063;
    wire N__47062;
    wire N__47061;
    wire N__47060;
    wire N__47059;
    wire N__47058;
    wire N__47057;
    wire N__47056;
    wire N__47055;
    wire N__47052;
    wire N__47047;
    wire N__47042;
    wire N__47033;
    wire N__47028;
    wire N__47021;
    wire N__47020;
    wire N__47015;
    wire N__47012;
    wire N__46997;
    wire N__46986;
    wire N__46979;
    wire N__46972;
    wire N__46959;
    wire N__46956;
    wire N__46951;
    wire N__46942;
    wire N__46939;
    wire N__46930;
    wire N__46929;
    wire N__46928;
    wire N__46927;
    wire N__46926;
    wire N__46925;
    wire N__46924;
    wire N__46923;
    wire N__46922;
    wire N__46919;
    wire N__46916;
    wire N__46905;
    wire N__46898;
    wire N__46891;
    wire N__46890;
    wire N__46887;
    wire N__46886;
    wire N__46885;
    wire N__46884;
    wire N__46881;
    wire N__46878;
    wire N__46875;
    wire N__46874;
    wire N__46871;
    wire N__46870;
    wire N__46867;
    wire N__46864;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46852;
    wire N__46849;
    wire N__46838;
    wire N__46831;
    wire N__46830;
    wire N__46829;
    wire N__46828;
    wire N__46827;
    wire N__46826;
    wire N__46825;
    wire N__46824;
    wire N__46823;
    wire N__46822;
    wire N__46819;
    wire N__46816;
    wire N__46813;
    wire N__46812;
    wire N__46811;
    wire N__46810;
    wire N__46807;
    wire N__46806;
    wire N__46805;
    wire N__46804;
    wire N__46803;
    wire N__46802;
    wire N__46801;
    wire N__46800;
    wire N__46799;
    wire N__46796;
    wire N__46795;
    wire N__46794;
    wire N__46791;
    wire N__46776;
    wire N__46773;
    wire N__46768;
    wire N__46765;
    wire N__46754;
    wire N__46751;
    wire N__46748;
    wire N__46747;
    wire N__46746;
    wire N__46745;
    wire N__46742;
    wire N__46735;
    wire N__46732;
    wire N__46729;
    wire N__46726;
    wire N__46719;
    wire N__46714;
    wire N__46709;
    wire N__46706;
    wire N__46699;
    wire N__46694;
    wire N__46687;
    wire N__46678;
    wire N__46675;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46665;
    wire N__46664;
    wire N__46663;
    wire N__46660;
    wire N__46657;
    wire N__46656;
    wire N__46653;
    wire N__46650;
    wire N__46647;
    wire N__46644;
    wire N__46643;
    wire N__46640;
    wire N__46635;
    wire N__46632;
    wire N__46629;
    wire N__46626;
    wire N__46623;
    wire N__46618;
    wire N__46615;
    wire N__46606;
    wire N__46603;
    wire N__46600;
    wire N__46599;
    wire N__46598;
    wire N__46595;
    wire N__46592;
    wire N__46589;
    wire N__46588;
    wire N__46587;
    wire N__46584;
    wire N__46581;
    wire N__46578;
    wire N__46575;
    wire N__46572;
    wire N__46569;
    wire N__46564;
    wire N__46555;
    wire N__46552;
    wire N__46549;
    wire N__46546;
    wire N__46545;
    wire N__46542;
    wire N__46539;
    wire N__46534;
    wire N__46533;
    wire N__46530;
    wire N__46527;
    wire N__46524;
    wire N__46521;
    wire N__46520;
    wire N__46517;
    wire N__46514;
    wire N__46511;
    wire N__46508;
    wire N__46501;
    wire N__46498;
    wire N__46495;
    wire N__46492;
    wire N__46489;
    wire N__46486;
    wire N__46483;
    wire N__46480;
    wire N__46477;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46462;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46435;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46420;
    wire N__46417;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46405;
    wire N__46402;
    wire N__46399;
    wire N__46396;
    wire N__46393;
    wire N__46390;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46357;
    wire N__46354;
    wire N__46351;
    wire N__46348;
    wire N__46345;
    wire N__46342;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46330;
    wire N__46327;
    wire N__46324;
    wire N__46321;
    wire N__46318;
    wire N__46315;
    wire N__46312;
    wire N__46309;
    wire N__46306;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46291;
    wire N__46288;
    wire N__46285;
    wire N__46282;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46245;
    wire N__46240;
    wire N__46237;
    wire N__46234;
    wire N__46233;
    wire N__46228;
    wire N__46225;
    wire N__46222;
    wire N__46221;
    wire N__46220;
    wire N__46219;
    wire N__46218;
    wire N__46215;
    wire N__46206;
    wire N__46201;
    wire N__46198;
    wire N__46197;
    wire N__46194;
    wire N__46191;
    wire N__46190;
    wire N__46187;
    wire N__46182;
    wire N__46181;
    wire N__46178;
    wire N__46175;
    wire N__46172;
    wire N__46169;
    wire N__46166;
    wire N__46159;
    wire N__46158;
    wire N__46153;
    wire N__46152;
    wire N__46151;
    wire N__46148;
    wire N__46143;
    wire N__46140;
    wire N__46135;
    wire N__46132;
    wire N__46129;
    wire N__46128;
    wire N__46127;
    wire N__46126;
    wire N__46125;
    wire N__46122;
    wire N__46113;
    wire N__46108;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46072;
    wire N__46069;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46051;
    wire N__46048;
    wire N__46047;
    wire N__46044;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46032;
    wire N__46027;
    wire N__46024;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46016;
    wire N__46015;
    wire N__46014;
    wire N__46013;
    wire N__46008;
    wire N__46005;
    wire N__46004;
    wire N__46001;
    wire N__46000;
    wire N__45997;
    wire N__45994;
    wire N__45991;
    wire N__45988;
    wire N__45985;
    wire N__45982;
    wire N__45979;
    wire N__45964;
    wire N__45961;
    wire N__45960;
    wire N__45959;
    wire N__45958;
    wire N__45955;
    wire N__45950;
    wire N__45947;
    wire N__45942;
    wire N__45937;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45929;
    wire N__45928;
    wire N__45927;
    wire N__45926;
    wire N__45923;
    wire N__45922;
    wire N__45919;
    wire N__45916;
    wire N__45915;
    wire N__45912;
    wire N__45911;
    wire N__45908;
    wire N__45907;
    wire N__45906;
    wire N__45905;
    wire N__45904;
    wire N__45903;
    wire N__45902;
    wire N__45899;
    wire N__45896;
    wire N__45893;
    wire N__45888;
    wire N__45881;
    wire N__45878;
    wire N__45875;
    wire N__45874;
    wire N__45873;
    wire N__45872;
    wire N__45869;
    wire N__45868;
    wire N__45865;
    wire N__45862;
    wire N__45861;
    wire N__45860;
    wire N__45855;
    wire N__45848;
    wire N__45841;
    wire N__45830;
    wire N__45819;
    wire N__45808;
    wire N__45805;
    wire N__45802;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45790;
    wire N__45787;
    wire N__45786;
    wire N__45783;
    wire N__45780;
    wire N__45779;
    wire N__45774;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45762;
    wire N__45757;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45739;
    wire N__45736;
    wire N__45735;
    wire N__45732;
    wire N__45731;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45717;
    wire N__45714;
    wire N__45709;
    wire N__45706;
    wire N__45705;
    wire N__45702;
    wire N__45701;
    wire N__45694;
    wire N__45691;
    wire N__45686;
    wire N__45683;
    wire N__45680;
    wire N__45673;
    wire N__45672;
    wire N__45669;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45656;
    wire N__45655;
    wire N__45654;
    wire N__45649;
    wire N__45646;
    wire N__45641;
    wire N__45638;
    wire N__45631;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45615;
    wire N__45610;
    wire N__45609;
    wire N__45606;
    wire N__45603;
    wire N__45602;
    wire N__45599;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45589;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45579;
    wire N__45576;
    wire N__45573;
    wire N__45562;
    wire N__45561;
    wire N__45560;
    wire N__45557;
    wire N__45556;
    wire N__45553;
    wire N__45552;
    wire N__45551;
    wire N__45550;
    wire N__45549;
    wire N__45548;
    wire N__45547;
    wire N__45546;
    wire N__45545;
    wire N__45540;
    wire N__45537;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45524;
    wire N__45521;
    wire N__45518;
    wire N__45515;
    wire N__45514;
    wire N__45513;
    wire N__45512;
    wire N__45511;
    wire N__45508;
    wire N__45505;
    wire N__45502;
    wire N__45499;
    wire N__45496;
    wire N__45491;
    wire N__45486;
    wire N__45483;
    wire N__45478;
    wire N__45471;
    wire N__45470;
    wire N__45467;
    wire N__45466;
    wire N__45465;
    wire N__45464;
    wire N__45463;
    wire N__45462;
    wire N__45461;
    wire N__45460;
    wire N__45459;
    wire N__45458;
    wire N__45457;
    wire N__45456;
    wire N__45455;
    wire N__45450;
    wire N__45447;
    wire N__45436;
    wire N__45431;
    wire N__45428;
    wire N__45425;
    wire N__45420;
    wire N__45409;
    wire N__45398;
    wire N__45379;
    wire N__45376;
    wire N__45375;
    wire N__45374;
    wire N__45371;
    wire N__45370;
    wire N__45365;
    wire N__45364;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45354;
    wire N__45353;
    wire N__45352;
    wire N__45349;
    wire N__45348;
    wire N__45343;
    wire N__45340;
    wire N__45337;
    wire N__45336;
    wire N__45335;
    wire N__45334;
    wire N__45333;
    wire N__45332;
    wire N__45329;
    wire N__45326;
    wire N__45323;
    wire N__45320;
    wire N__45317;
    wire N__45316;
    wire N__45315;
    wire N__45314;
    wire N__45313;
    wire N__45312;
    wire N__45311;
    wire N__45306;
    wire N__45303;
    wire N__45300;
    wire N__45297;
    wire N__45294;
    wire N__45291;
    wire N__45290;
    wire N__45287;
    wire N__45284;
    wire N__45281;
    wire N__45276;
    wire N__45271;
    wire N__45268;
    wire N__45265;
    wire N__45260;
    wire N__45257;
    wire N__45252;
    wire N__45249;
    wire N__45246;
    wire N__45243;
    wire N__45240;
    wire N__45223;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45199;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45169;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45151;
    wire N__45148;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45097;
    wire N__45096;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45064;
    wire N__45061;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45046;
    wire N__45043;
    wire N__45040;
    wire N__45037;
    wire N__45034;
    wire N__45031;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45013;
    wire N__45010;
    wire N__45007;
    wire N__45006;
    wire N__45003;
    wire N__45000;
    wire N__44995;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44987;
    wire N__44984;
    wire N__44981;
    wire N__44978;
    wire N__44975;
    wire N__44972;
    wire N__44971;
    wire N__44968;
    wire N__44963;
    wire N__44960;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44944;
    wire N__44941;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44933;
    wire N__44930;
    wire N__44927;
    wire N__44924;
    wire N__44919;
    wire N__44914;
    wire N__44911;
    wire N__44908;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44898;
    wire N__44895;
    wire N__44890;
    wire N__44887;
    wire N__44884;
    wire N__44883;
    wire N__44880;
    wire N__44877;
    wire N__44876;
    wire N__44873;
    wire N__44870;
    wire N__44867;
    wire N__44862;
    wire N__44857;
    wire N__44854;
    wire N__44853;
    wire N__44850;
    wire N__44847;
    wire N__44844;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44823;
    wire N__44820;
    wire N__44817;
    wire N__44814;
    wire N__44809;
    wire N__44806;
    wire N__44805;
    wire N__44804;
    wire N__44801;
    wire N__44798;
    wire N__44795;
    wire N__44790;
    wire N__44785;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44766;
    wire N__44761;
    wire N__44758;
    wire N__44757;
    wire N__44756;
    wire N__44753;
    wire N__44748;
    wire N__44743;
    wire N__44740;
    wire N__44737;
    wire N__44736;
    wire N__44733;
    wire N__44730;
    wire N__44727;
    wire N__44722;
    wire N__44721;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44704;
    wire N__44701;
    wire N__44698;
    wire N__44695;
    wire N__44694;
    wire N__44693;
    wire N__44692;
    wire N__44687;
    wire N__44684;
    wire N__44681;
    wire N__44680;
    wire N__44677;
    wire N__44674;
    wire N__44671;
    wire N__44668;
    wire N__44665;
    wire N__44664;
    wire N__44657;
    wire N__44654;
    wire N__44651;
    wire N__44648;
    wire N__44641;
    wire N__44640;
    wire N__44637;
    wire N__44634;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44624;
    wire N__44619;
    wire N__44618;
    wire N__44615;
    wire N__44612;
    wire N__44609;
    wire N__44602;
    wire N__44601;
    wire N__44598;
    wire N__44597;
    wire N__44594;
    wire N__44591;
    wire N__44588;
    wire N__44585;
    wire N__44582;
    wire N__44579;
    wire N__44576;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44562;
    wire N__44557;
    wire N__44554;
    wire N__44553;
    wire N__44552;
    wire N__44549;
    wire N__44546;
    wire N__44543;
    wire N__44542;
    wire N__44541;
    wire N__44536;
    wire N__44533;
    wire N__44532;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44512;
    wire N__44503;
    wire N__44500;
    wire N__44497;
    wire N__44494;
    wire N__44491;
    wire N__44490;
    wire N__44487;
    wire N__44484;
    wire N__44479;
    wire N__44476;
    wire N__44475;
    wire N__44472;
    wire N__44469;
    wire N__44466;
    wire N__44463;
    wire N__44462;
    wire N__44457;
    wire N__44454;
    wire N__44451;
    wire N__44446;
    wire N__44443;
    wire N__44440;
    wire N__44437;
    wire N__44436;
    wire N__44435;
    wire N__44432;
    wire N__44429;
    wire N__44426;
    wire N__44421;
    wire N__44416;
    wire N__44413;
    wire N__44410;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44398;
    wire N__44395;
    wire N__44394;
    wire N__44393;
    wire N__44388;
    wire N__44385;
    wire N__44382;
    wire N__44377;
    wire N__44374;
    wire N__44371;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44359;
    wire N__44356;
    wire N__44355;
    wire N__44354;
    wire N__44349;
    wire N__44346;
    wire N__44343;
    wire N__44338;
    wire N__44335;
    wire N__44332;
    wire N__44331;
    wire N__44328;
    wire N__44325;
    wire N__44320;
    wire N__44317;
    wire N__44316;
    wire N__44313;
    wire N__44310;
    wire N__44309;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44293;
    wire N__44290;
    wire N__44289;
    wire N__44286;
    wire N__44283;
    wire N__44278;
    wire N__44275;
    wire N__44272;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44264;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44248;
    wire N__44245;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44233;
    wire N__44230;
    wire N__44227;
    wire N__44226;
    wire N__44221;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44185;
    wire N__44182;
    wire N__44181;
    wire N__44176;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44161;
    wire N__44158;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44142;
    wire N__44139;
    wire N__44134;
    wire N__44131;
    wire N__44128;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44120;
    wire N__44117;
    wire N__44114;
    wire N__44111;
    wire N__44106;
    wire N__44101;
    wire N__44098;
    wire N__44095;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44083;
    wire N__44080;
    wire N__44079;
    wire N__44076;
    wire N__44073;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44058;
    wire N__44053;
    wire N__44050;
    wire N__44047;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44035;
    wire N__44032;
    wire N__44031;
    wire N__44026;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44011;
    wire N__44008;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43973;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43957;
    wire N__43954;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43946;
    wire N__43941;
    wire N__43938;
    wire N__43935;
    wire N__43930;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43916;
    wire N__43911;
    wire N__43908;
    wire N__43903;
    wire N__43900;
    wire N__43899;
    wire N__43898;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43882;
    wire N__43879;
    wire N__43878;
    wire N__43873;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43863;
    wire N__43858;
    wire N__43855;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43843;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43833;
    wire N__43828;
    wire N__43825;
    wire N__43824;
    wire N__43823;
    wire N__43822;
    wire N__43821;
    wire N__43820;
    wire N__43819;
    wire N__43818;
    wire N__43817;
    wire N__43816;
    wire N__43815;
    wire N__43814;
    wire N__43813;
    wire N__43812;
    wire N__43811;
    wire N__43810;
    wire N__43809;
    wire N__43808;
    wire N__43799;
    wire N__43790;
    wire N__43781;
    wire N__43780;
    wire N__43779;
    wire N__43778;
    wire N__43777;
    wire N__43776;
    wire N__43775;
    wire N__43774;
    wire N__43773;
    wire N__43772;
    wire N__43771;
    wire N__43770;
    wire N__43769;
    wire N__43764;
    wire N__43755;
    wire N__43748;
    wire N__43739;
    wire N__43730;
    wire N__43721;
    wire N__43718;
    wire N__43715;
    wire N__43710;
    wire N__43705;
    wire N__43700;
    wire N__43697;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43676;
    wire N__43675;
    wire N__43670;
    wire N__43667;
    wire N__43664;
    wire N__43661;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43649;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43637;
    wire N__43630;
    wire N__43627;
    wire N__43626;
    wire N__43621;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43606;
    wire N__43603;
    wire N__43602;
    wire N__43597;
    wire N__43596;
    wire N__43593;
    wire N__43590;
    wire N__43587;
    wire N__43582;
    wire N__43579;
    wire N__43578;
    wire N__43575;
    wire N__43572;
    wire N__43571;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43555;
    wire N__43552;
    wire N__43551;
    wire N__43548;
    wire N__43545;
    wire N__43544;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43528;
    wire N__43525;
    wire N__43524;
    wire N__43519;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43504;
    wire N__43501;
    wire N__43500;
    wire N__43495;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43485;
    wire N__43480;
    wire N__43477;
    wire N__43476;
    wire N__43473;
    wire N__43470;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43411;
    wire N__43408;
    wire N__43405;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43393;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43377;
    wire N__43376;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43366;
    wire N__43363;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43345;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43335;
    wire N__43332;
    wire N__43329;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43308;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43298;
    wire N__43297;
    wire N__43292;
    wire N__43289;
    wire N__43286;
    wire N__43281;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43264;
    wire N__43263;
    wire N__43260;
    wire N__43259;
    wire N__43256;
    wire N__43253;
    wire N__43250;
    wire N__43249;
    wire N__43244;
    wire N__43239;
    wire N__43234;
    wire N__43231;
    wire N__43228;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43208;
    wire N__43203;
    wire N__43200;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43150;
    wire N__43149;
    wire N__43148;
    wire N__43145;
    wire N__43144;
    wire N__43143;
    wire N__43142;
    wire N__43141;
    wire N__43140;
    wire N__43139;
    wire N__43138;
    wire N__43137;
    wire N__43136;
    wire N__43135;
    wire N__43134;
    wire N__43133;
    wire N__43132;
    wire N__43131;
    wire N__43130;
    wire N__43129;
    wire N__43128;
    wire N__43127;
    wire N__43126;
    wire N__43125;
    wire N__43124;
    wire N__43123;
    wire N__43122;
    wire N__43121;
    wire N__43118;
    wire N__43115;
    wire N__43112;
    wire N__43109;
    wire N__43106;
    wire N__43097;
    wire N__43096;
    wire N__43095;
    wire N__43094;
    wire N__43093;
    wire N__43092;
    wire N__43091;
    wire N__43090;
    wire N__43089;
    wire N__43082;
    wire N__43073;
    wire N__43064;
    wire N__43055;
    wire N__43048;
    wire N__43043;
    wire N__43042;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43022;
    wire N__43013;
    wire N__43006;
    wire N__43001;
    wire N__42998;
    wire N__42995;
    wire N__42992;
    wire N__42979;
    wire N__42970;
    wire N__42967;
    wire N__42964;
    wire N__42963;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42955;
    wire N__42954;
    wire N__42951;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42931;
    wire N__42928;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42918;
    wire N__42913;
    wire N__42910;
    wire N__42909;
    wire N__42906;
    wire N__42903;
    wire N__42898;
    wire N__42895;
    wire N__42894;
    wire N__42891;
    wire N__42888;
    wire N__42885;
    wire N__42882;
    wire N__42879;
    wire N__42874;
    wire N__42871;
    wire N__42870;
    wire N__42867;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42850;
    wire N__42847;
    wire N__42846;
    wire N__42843;
    wire N__42842;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42827;
    wire N__42820;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42808;
    wire N__42805;
    wire N__42802;
    wire N__42801;
    wire N__42796;
    wire N__42793;
    wire N__42790;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42778;
    wire N__42775;
    wire N__42774;
    wire N__42773;
    wire N__42770;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42757;
    wire N__42752;
    wire N__42749;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42727;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42717;
    wire N__42712;
    wire N__42709;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42699;
    wire N__42694;
    wire N__42691;
    wire N__42690;
    wire N__42685;
    wire N__42682;
    wire N__42681;
    wire N__42676;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42661;
    wire N__42658;
    wire N__42655;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42645;
    wire N__42644;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42631;
    wire N__42628;
    wire N__42619;
    wire N__42618;
    wire N__42613;
    wire N__42610;
    wire N__42609;
    wire N__42606;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42592;
    wire N__42591;
    wire N__42588;
    wire N__42583;
    wire N__42580;
    wire N__42577;
    wire N__42574;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42562;
    wire N__42559;
    wire N__42556;
    wire N__42555;
    wire N__42550;
    wire N__42547;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42526;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42508;
    wire N__42505;
    wire N__42502;
    wire N__42499;
    wire N__42496;
    wire N__42495;
    wire N__42490;
    wire N__42487;
    wire N__42486;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42460;
    wire N__42457;
    wire N__42454;
    wire N__42451;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42439;
    wire N__42436;
    wire N__42433;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42421;
    wire N__42418;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42406;
    wire N__42403;
    wire N__42400;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42382;
    wire N__42379;
    wire N__42378;
    wire N__42375;
    wire N__42372;
    wire N__42367;
    wire N__42364;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42352;
    wire N__42349;
    wire N__42346;
    wire N__42345;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42328;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42313;
    wire N__42310;
    wire N__42307;
    wire N__42306;
    wire N__42303;
    wire N__42302;
    wire N__42299;
    wire N__42296;
    wire N__42293;
    wire N__42286;
    wire N__42285;
    wire N__42284;
    wire N__42283;
    wire N__42282;
    wire N__42281;
    wire N__42280;
    wire N__42279;
    wire N__42276;
    wire N__42273;
    wire N__42272;
    wire N__42271;
    wire N__42268;
    wire N__42267;
    wire N__42256;
    wire N__42253;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42239;
    wire N__42228;
    wire N__42223;
    wire N__42220;
    wire N__42217;
    wire N__42216;
    wire N__42215;
    wire N__42214;
    wire N__42213;
    wire N__42212;
    wire N__42209;
    wire N__42206;
    wire N__42205;
    wire N__42204;
    wire N__42203;
    wire N__42202;
    wire N__42201;
    wire N__42200;
    wire N__42197;
    wire N__42194;
    wire N__42193;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42181;
    wire N__42178;
    wire N__42173;
    wire N__42162;
    wire N__42157;
    wire N__42154;
    wire N__42149;
    wire N__42136;
    wire N__42135;
    wire N__42132;
    wire N__42129;
    wire N__42124;
    wire N__42121;
    wire N__42118;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42106;
    wire N__42103;
    wire N__42100;
    wire N__42097;
    wire N__42094;
    wire N__42091;
    wire N__42088;
    wire N__42085;
    wire N__42082;
    wire N__42079;
    wire N__42076;
    wire N__42073;
    wire N__42070;
    wire N__42067;
    wire N__42064;
    wire N__42061;
    wire N__42058;
    wire N__42055;
    wire N__42052;
    wire N__42049;
    wire N__42046;
    wire N__42045;
    wire N__42042;
    wire N__42039;
    wire N__42034;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42016;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42006;
    wire N__42003;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41989;
    wire N__41986;
    wire N__41983;
    wire N__41980;
    wire N__41977;
    wire N__41974;
    wire N__41971;
    wire N__41968;
    wire N__41967;
    wire N__41964;
    wire N__41963;
    wire N__41960;
    wire N__41957;
    wire N__41956;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41941;
    wire N__41932;
    wire N__41931;
    wire N__41926;
    wire N__41923;
    wire N__41922;
    wire N__41919;
    wire N__41918;
    wire N__41915;
    wire N__41912;
    wire N__41911;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41887;
    wire N__41884;
    wire N__41883;
    wire N__41878;
    wire N__41875;
    wire N__41874;
    wire N__41869;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41861;
    wire N__41860;
    wire N__41857;
    wire N__41854;
    wire N__41851;
    wire N__41848;
    wire N__41839;
    wire N__41836;
    wire N__41833;
    wire N__41830;
    wire N__41827;
    wire N__41824;
    wire N__41823;
    wire N__41818;
    wire N__41815;
    wire N__41812;
    wire N__41809;
    wire N__41808;
    wire N__41807;
    wire N__41806;
    wire N__41805;
    wire N__41804;
    wire N__41803;
    wire N__41802;
    wire N__41801;
    wire N__41800;
    wire N__41799;
    wire N__41798;
    wire N__41787;
    wire N__41782;
    wire N__41781;
    wire N__41780;
    wire N__41779;
    wire N__41778;
    wire N__41777;
    wire N__41776;
    wire N__41775;
    wire N__41774;
    wire N__41773;
    wire N__41772;
    wire N__41771;
    wire N__41770;
    wire N__41769;
    wire N__41768;
    wire N__41765;
    wire N__41764;
    wire N__41763;
    wire N__41762;
    wire N__41761;
    wire N__41752;
    wire N__41751;
    wire N__41750;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41732;
    wire N__41719;
    wire N__41716;
    wire N__41707;
    wire N__41700;
    wire N__41699;
    wire N__41698;
    wire N__41695;
    wire N__41688;
    wire N__41681;
    wire N__41672;
    wire N__41667;
    wire N__41656;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41648;
    wire N__41647;
    wire N__41638;
    wire N__41637;
    wire N__41636;
    wire N__41635;
    wire N__41634;
    wire N__41633;
    wire N__41632;
    wire N__41631;
    wire N__41630;
    wire N__41629;
    wire N__41628;
    wire N__41627;
    wire N__41626;
    wire N__41625;
    wire N__41624;
    wire N__41623;
    wire N__41622;
    wire N__41621;
    wire N__41618;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41600;
    wire N__41597;
    wire N__41596;
    wire N__41595;
    wire N__41594;
    wire N__41593;
    wire N__41586;
    wire N__41583;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41568;
    wire N__41565;
    wire N__41562;
    wire N__41555;
    wire N__41546;
    wire N__41543;
    wire N__41538;
    wire N__41535;
    wire N__41526;
    wire N__41521;
    wire N__41510;
    wire N__41503;
    wire N__41502;
    wire N__41499;
    wire N__41498;
    wire N__41495;
    wire N__41492;
    wire N__41489;
    wire N__41488;
    wire N__41485;
    wire N__41482;
    wire N__41479;
    wire N__41476;
    wire N__41467;
    wire N__41466;
    wire N__41461;
    wire N__41458;
    wire N__41455;
    wire N__41452;
    wire N__41449;
    wire N__41448;
    wire N__41445;
    wire N__41444;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41434;
    wire N__41433;
    wire N__41432;
    wire N__41429;
    wire N__41426;
    wire N__41421;
    wire N__41418;
    wire N__41415;
    wire N__41412;
    wire N__41409;
    wire N__41402;
    wire N__41395;
    wire N__41392;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41380;
    wire N__41377;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41365;
    wire N__41364;
    wire N__41363;
    wire N__41362;
    wire N__41361;
    wire N__41360;
    wire N__41359;
    wire N__41358;
    wire N__41355;
    wire N__41348;
    wire N__41339;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41320;
    wire N__41319;
    wire N__41318;
    wire N__41317;
    wire N__41312;
    wire N__41311;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41296;
    wire N__41291;
    wire N__41286;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41263;
    wire N__41262;
    wire N__41261;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41246;
    wire N__41243;
    wire N__41240;
    wire N__41237;
    wire N__41234;
    wire N__41227;
    wire N__41224;
    wire N__41223;
    wire N__41222;
    wire N__41219;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41200;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41190;
    wire N__41189;
    wire N__41186;
    wire N__41181;
    wire N__41176;
    wire N__41173;
    wire N__41170;
    wire N__41169;
    wire N__41168;
    wire N__41165;
    wire N__41160;
    wire N__41155;
    wire N__41152;
    wire N__41149;
    wire N__41146;
    wire N__41143;
    wire N__41140;
    wire N__41139;
    wire N__41138;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41125;
    wire N__41122;
    wire N__41117;
    wire N__41114;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41100;
    wire N__41097;
    wire N__41096;
    wire N__41093;
    wire N__41090;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41077;
    wire N__41068;
    wire N__41065;
    wire N__41062;
    wire N__41061;
    wire N__41060;
    wire N__41057;
    wire N__41056;
    wire N__41055;
    wire N__41054;
    wire N__41051;
    wire N__41050;
    wire N__41049;
    wire N__41046;
    wire N__41045;
    wire N__41044;
    wire N__41043;
    wire N__41042;
    wire N__41041;
    wire N__41040;
    wire N__41039;
    wire N__41036;
    wire N__41035;
    wire N__41034;
    wire N__41033;
    wire N__41032;
    wire N__41031;
    wire N__41030;
    wire N__41029;
    wire N__41026;
    wire N__41025;
    wire N__41024;
    wire N__41023;
    wire N__41022;
    wire N__41019;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40987;
    wire N__40984;
    wire N__40975;
    wire N__40974;
    wire N__40973;
    wire N__40972;
    wire N__40969;
    wire N__40966;
    wire N__40963;
    wire N__40960;
    wire N__40951;
    wire N__40946;
    wire N__40943;
    wire N__40938;
    wire N__40929;
    wire N__40924;
    wire N__40917;
    wire N__40910;
    wire N__40891;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40867;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40857;
    wire N__40856;
    wire N__40853;
    wire N__40848;
    wire N__40843;
    wire N__40840;
    wire N__40839;
    wire N__40836;
    wire N__40835;
    wire N__40832;
    wire N__40827;
    wire N__40822;
    wire N__40821;
    wire N__40820;
    wire N__40819;
    wire N__40818;
    wire N__40817;
    wire N__40816;
    wire N__40815;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40788;
    wire N__40787;
    wire N__40786;
    wire N__40785;
    wire N__40784;
    wire N__40783;
    wire N__40782;
    wire N__40781;
    wire N__40780;
    wire N__40779;
    wire N__40778;
    wire N__40777;
    wire N__40776;
    wire N__40771;
    wire N__40768;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40750;
    wire N__40745;
    wire N__40740;
    wire N__40733;
    wire N__40726;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40685;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40675;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40663;
    wire N__40660;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40638;
    wire N__40635;
    wire N__40634;
    wire N__40631;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40613;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40584;
    wire N__40581;
    wire N__40578;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40563;
    wire N__40560;
    wire N__40557;
    wire N__40552;
    wire N__40551;
    wire N__40550;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40534;
    wire N__40531;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40523;
    wire N__40518;
    wire N__40515;
    wire N__40512;
    wire N__40507;
    wire N__40504;
    wire N__40501;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40491;
    wire N__40486;
    wire N__40483;
    wire N__40482;
    wire N__40481;
    wire N__40480;
    wire N__40479;
    wire N__40478;
    wire N__40477;
    wire N__40476;
    wire N__40467;
    wire N__40466;
    wire N__40465;
    wire N__40464;
    wire N__40463;
    wire N__40462;
    wire N__40461;
    wire N__40460;
    wire N__40459;
    wire N__40458;
    wire N__40457;
    wire N__40456;
    wire N__40455;
    wire N__40454;
    wire N__40453;
    wire N__40444;
    wire N__40443;
    wire N__40442;
    wire N__40441;
    wire N__40440;
    wire N__40437;
    wire N__40432;
    wire N__40423;
    wire N__40414;
    wire N__40405;
    wire N__40404;
    wire N__40403;
    wire N__40402;
    wire N__40401;
    wire N__40398;
    wire N__40389;
    wire N__40382;
    wire N__40379;
    wire N__40376;
    wire N__40367;
    wire N__40358;
    wire N__40353;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40327;
    wire N__40326;
    wire N__40325;
    wire N__40322;
    wire N__40319;
    wire N__40318;
    wire N__40315;
    wire N__40310;
    wire N__40307;
    wire N__40304;
    wire N__40301;
    wire N__40298;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40279;
    wire N__40278;
    wire N__40275;
    wire N__40272;
    wire N__40267;
    wire N__40264;
    wire N__40263;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40239;
    wire N__40238;
    wire N__40235;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40216;
    wire N__40213;
    wire N__40210;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40202;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40186;
    wire N__40183;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40175;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40159;
    wire N__40156;
    wire N__40155;
    wire N__40154;
    wire N__40149;
    wire N__40146;
    wire N__40143;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40131;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40116;
    wire N__40111;
    wire N__40108;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40096;
    wire N__40095;
    wire N__40092;
    wire N__40089;
    wire N__40086;
    wire N__40081;
    wire N__40078;
    wire N__40077;
    wire N__40076;
    wire N__40071;
    wire N__40068;
    wire N__40065;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40051;
    wire N__40050;
    wire N__40049;
    wire N__40046;
    wire N__40043;
    wire N__40040;
    wire N__40037;
    wire N__40034;
    wire N__40027;
    wire N__40024;
    wire N__40023;
    wire N__40020;
    wire N__40017;
    wire N__40016;
    wire N__40013;
    wire N__40010;
    wire N__40007;
    wire N__40004;
    wire N__40001;
    wire N__39994;
    wire N__39991;
    wire N__39988;
    wire N__39987;
    wire N__39984;
    wire N__39981;
    wire N__39980;
    wire N__39975;
    wire N__39972;
    wire N__39969;
    wire N__39964;
    wire N__39961;
    wire N__39960;
    wire N__39955;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39940;
    wire N__39937;
    wire N__39936;
    wire N__39931;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39916;
    wire N__39913;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39901;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39886;
    wire N__39883;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39871;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39842;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39826;
    wire N__39823;
    wire N__39820;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39812;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39768;
    wire N__39763;
    wire N__39760;
    wire N__39759;
    wire N__39756;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39746;
    wire N__39743;
    wire N__39740;
    wire N__39737;
    wire N__39734;
    wire N__39727;
    wire N__39724;
    wire N__39723;
    wire N__39722;
    wire N__39717;
    wire N__39714;
    wire N__39711;
    wire N__39706;
    wire N__39703;
    wire N__39702;
    wire N__39697;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39682;
    wire N__39679;
    wire N__39678;
    wire N__39675;
    wire N__39674;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39660;
    wire N__39655;
    wire N__39652;
    wire N__39651;
    wire N__39648;
    wire N__39645;
    wire N__39640;
    wire N__39639;
    wire N__39636;
    wire N__39633;
    wire N__39630;
    wire N__39625;
    wire N__39622;
    wire N__39621;
    wire N__39618;
    wire N__39615;
    wire N__39610;
    wire N__39609;
    wire N__39606;
    wire N__39603;
    wire N__39600;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39581;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39565;
    wire N__39562;
    wire N__39559;
    wire N__39556;
    wire N__39555;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39545;
    wire N__39542;
    wire N__39539;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39490;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39450;
    wire N__39449;
    wire N__39448;
    wire N__39447;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39424;
    wire N__39423;
    wire N__39422;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39391;
    wire N__39388;
    wire N__39385;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39373;
    wire N__39372;
    wire N__39367;
    wire N__39364;
    wire N__39361;
    wire N__39358;
    wire N__39357;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39340;
    wire N__39339;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39313;
    wire N__39310;
    wire N__39307;
    wire N__39304;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39296;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39284;
    wire N__39281;
    wire N__39278;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39262;
    wire N__39259;
    wire N__39258;
    wire N__39253;
    wire N__39250;
    wire N__39249;
    wire N__39244;
    wire N__39241;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39229;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39205;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39193;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39165;
    wire N__39162;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39082;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39025;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38910;
    wire N__38909;
    wire N__38904;
    wire N__38901;
    wire N__38896;
    wire N__38895;
    wire N__38892;
    wire N__38889;
    wire N__38884;
    wire N__38881;
    wire N__38878;
    wire N__38875;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38863;
    wire N__38860;
    wire N__38857;
    wire N__38856;
    wire N__38855;
    wire N__38852;
    wire N__38851;
    wire N__38850;
    wire N__38849;
    wire N__38846;
    wire N__38845;
    wire N__38844;
    wire N__38843;
    wire N__38840;
    wire N__38839;
    wire N__38838;
    wire N__38837;
    wire N__38834;
    wire N__38829;
    wire N__38824;
    wire N__38819;
    wire N__38808;
    wire N__38805;
    wire N__38794;
    wire N__38793;
    wire N__38792;
    wire N__38791;
    wire N__38790;
    wire N__38783;
    wire N__38782;
    wire N__38781;
    wire N__38780;
    wire N__38777;
    wire N__38776;
    wire N__38773;
    wire N__38772;
    wire N__38771;
    wire N__38770;
    wire N__38769;
    wire N__38768;
    wire N__38765;
    wire N__38760;
    wire N__38757;
    wire N__38752;
    wire N__38747;
    wire N__38738;
    wire N__38735;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38695;
    wire N__38692;
    wire N__38689;
    wire N__38688;
    wire N__38685;
    wire N__38684;
    wire N__38683;
    wire N__38680;
    wire N__38677;
    wire N__38674;
    wire N__38671;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38644;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38626;
    wire N__38623;
    wire N__38622;
    wire N__38621;
    wire N__38616;
    wire N__38613;
    wire N__38608;
    wire N__38607;
    wire N__38606;
    wire N__38603;
    wire N__38598;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38572;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38564;
    wire N__38561;
    wire N__38558;
    wire N__38555;
    wire N__38548;
    wire N__38547;
    wire N__38546;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38536;
    wire N__38533;
    wire N__38524;
    wire N__38523;
    wire N__38522;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38512;
    wire N__38509;
    wire N__38500;
    wire N__38499;
    wire N__38496;
    wire N__38495;
    wire N__38494;
    wire N__38491;
    wire N__38488;
    wire N__38485;
    wire N__38482;
    wire N__38473;
    wire N__38472;
    wire N__38471;
    wire N__38470;
    wire N__38469;
    wire N__38468;
    wire N__38467;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38448;
    wire N__38445;
    wire N__38434;
    wire N__38431;
    wire N__38430;
    wire N__38429;
    wire N__38428;
    wire N__38427;
    wire N__38426;
    wire N__38423;
    wire N__38420;
    wire N__38419;
    wire N__38418;
    wire N__38417;
    wire N__38416;
    wire N__38415;
    wire N__38414;
    wire N__38411;
    wire N__38400;
    wire N__38387;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38364;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38352;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38332;
    wire N__38331;
    wire N__38326;
    wire N__38323;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38312;
    wire N__38309;
    wire N__38306;
    wire N__38303;
    wire N__38296;
    wire N__38295;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38279;
    wire N__38274;
    wire N__38271;
    wire N__38266;
    wire N__38263;
    wire N__38260;
    wire N__38259;
    wire N__38258;
    wire N__38257;
    wire N__38256;
    wire N__38255;
    wire N__38254;
    wire N__38247;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38237;
    wire N__38234;
    wire N__38231;
    wire N__38228;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38202;
    wire N__38199;
    wire N__38196;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38178;
    wire N__38175;
    wire N__38174;
    wire N__38171;
    wire N__38168;
    wire N__38165;
    wire N__38162;
    wire N__38159;
    wire N__38156;
    wire N__38155;
    wire N__38154;
    wire N__38151;
    wire N__38146;
    wire N__38141;
    wire N__38138;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38103;
    wire N__38100;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38090;
    wire N__38087;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38069;
    wire N__38064;
    wire N__38059;
    wire N__38058;
    wire N__38057;
    wire N__38054;
    wire N__38051;
    wire N__38048;
    wire N__38041;
    wire N__38038;
    wire N__38037;
    wire N__38036;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38004;
    wire N__38001;
    wire N__37994;
    wire N__37991;
    wire N__37984;
    wire N__37983;
    wire N__37980;
    wire N__37979;
    wire N__37978;
    wire N__37977;
    wire N__37976;
    wire N__37975;
    wire N__37974;
    wire N__37973;
    wire N__37972;
    wire N__37971;
    wire N__37970;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37954;
    wire N__37951;
    wire N__37950;
    wire N__37949;
    wire N__37948;
    wire N__37947;
    wire N__37946;
    wire N__37945;
    wire N__37944;
    wire N__37943;
    wire N__37942;
    wire N__37941;
    wire N__37940;
    wire N__37939;
    wire N__37938;
    wire N__37937;
    wire N__37936;
    wire N__37935;
    wire N__37934;
    wire N__37933;
    wire N__37932;
    wire N__37919;
    wire N__37916;
    wire N__37911;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37893;
    wire N__37892;
    wire N__37889;
    wire N__37888;
    wire N__37885;
    wire N__37884;
    wire N__37883;
    wire N__37882;
    wire N__37879;
    wire N__37878;
    wire N__37877;
    wire N__37874;
    wire N__37873;
    wire N__37872;
    wire N__37871;
    wire N__37868;
    wire N__37867;
    wire N__37860;
    wire N__37851;
    wire N__37848;
    wire N__37839;
    wire N__37838;
    wire N__37837;
    wire N__37834;
    wire N__37833;
    wire N__37828;
    wire N__37817;
    wire N__37806;
    wire N__37793;
    wire N__37792;
    wire N__37791;
    wire N__37786;
    wire N__37781;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37761;
    wire N__37756;
    wire N__37751;
    wire N__37738;
    wire N__37735;
    wire N__37732;
    wire N__37729;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37714;
    wire N__37713;
    wire N__37710;
    wire N__37709;
    wire N__37708;
    wire N__37707;
    wire N__37706;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37694;
    wire N__37693;
    wire N__37692;
    wire N__37689;
    wire N__37688;
    wire N__37687;
    wire N__37686;
    wire N__37683;
    wire N__37682;
    wire N__37681;
    wire N__37674;
    wire N__37673;
    wire N__37672;
    wire N__37671;
    wire N__37670;
    wire N__37669;
    wire N__37668;
    wire N__37667;
    wire N__37666;
    wire N__37665;
    wire N__37664;
    wire N__37663;
    wire N__37660;
    wire N__37655;
    wire N__37652;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37631;
    wire N__37630;
    wire N__37629;
    wire N__37628;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37618;
    wire N__37615;
    wire N__37614;
    wire N__37613;
    wire N__37612;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37588;
    wire N__37583;
    wire N__37578;
    wire N__37573;
    wire N__37556;
    wire N__37545;
    wire N__37542;
    wire N__37537;
    wire N__37530;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37514;
    wire N__37501;
    wire N__37500;
    wire N__37499;
    wire N__37498;
    wire N__37497;
    wire N__37496;
    wire N__37495;
    wire N__37494;
    wire N__37493;
    wire N__37492;
    wire N__37489;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37475;
    wire N__37464;
    wire N__37461;
    wire N__37460;
    wire N__37457;
    wire N__37456;
    wire N__37455;
    wire N__37454;
    wire N__37453;
    wire N__37452;
    wire N__37451;
    wire N__37450;
    wire N__37449;
    wire N__37448;
    wire N__37447;
    wire N__37446;
    wire N__37445;
    wire N__37444;
    wire N__37443;
    wire N__37442;
    wire N__37441;
    wire N__37440;
    wire N__37439;
    wire N__37438;
    wire N__37435;
    wire N__37432;
    wire N__37427;
    wire N__37424;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37404;
    wire N__37387;
    wire N__37384;
    wire N__37377;
    wire N__37372;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37351;
    wire N__37344;
    wire N__37327;
    wire N__37326;
    wire N__37325;
    wire N__37324;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37316;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37308;
    wire N__37307;
    wire N__37304;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37290;
    wire N__37289;
    wire N__37288;
    wire N__37287;
    wire N__37286;
    wire N__37285;
    wire N__37284;
    wire N__37283;
    wire N__37282;
    wire N__37277;
    wire N__37274;
    wire N__37273;
    wire N__37272;
    wire N__37271;
    wire N__37270;
    wire N__37269;
    wire N__37268;
    wire N__37267;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37246;
    wire N__37235;
    wire N__37234;
    wire N__37233;
    wire N__37232;
    wire N__37231;
    wire N__37230;
    wire N__37227;
    wire N__37224;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37196;
    wire N__37191;
    wire N__37188;
    wire N__37183;
    wire N__37178;
    wire N__37175;
    wire N__37166;
    wire N__37161;
    wire N__37158;
    wire N__37151;
    wire N__37148;
    wire N__37143;
    wire N__37140;
    wire N__37123;
    wire N__37120;
    wire N__37117;
    wire N__37114;
    wire N__37111;
    wire N__37108;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37100;
    wire N__37095;
    wire N__37092;
    wire N__37091;
    wire N__37086;
    wire N__37083;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37073;
    wire N__37070;
    wire N__37067;
    wire N__37060;
    wire N__37057;
    wire N__37054;
    wire N__37051;
    wire N__37050;
    wire N__37047;
    wire N__37044;
    wire N__37043;
    wire N__37042;
    wire N__37037;
    wire N__37034;
    wire N__37031;
    wire N__37026;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37014;
    wire N__37011;
    wire N__37008;
    wire N__37005;
    wire N__37000;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36976;
    wire N__36973;
    wire N__36972;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36958;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36934;
    wire N__36931;
    wire N__36930;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36916;
    wire N__36915;
    wire N__36912;
    wire N__36909;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36891;
    wire N__36888;
    wire N__36885;
    wire N__36880;
    wire N__36879;
    wire N__36876;
    wire N__36873;
    wire N__36870;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36835;
    wire N__36834;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36820;
    wire N__36817;
    wire N__36814;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36799;
    wire N__36796;
    wire N__36795;
    wire N__36792;
    wire N__36789;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36766;
    wire N__36763;
    wire N__36762;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36754;
    wire N__36751;
    wire N__36750;
    wire N__36749;
    wire N__36748;
    wire N__36747;
    wire N__36746;
    wire N__36745;
    wire N__36744;
    wire N__36743;
    wire N__36740;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36730;
    wire N__36729;
    wire N__36728;
    wire N__36727;
    wire N__36726;
    wire N__36725;
    wire N__36724;
    wire N__36723;
    wire N__36722;
    wire N__36721;
    wire N__36720;
    wire N__36719;
    wire N__36716;
    wire N__36709;
    wire N__36700;
    wire N__36699;
    wire N__36698;
    wire N__36697;
    wire N__36696;
    wire N__36695;
    wire N__36694;
    wire N__36693;
    wire N__36692;
    wire N__36691;
    wire N__36690;
    wire N__36689;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36677;
    wire N__36674;
    wire N__36665;
    wire N__36656;
    wire N__36649;
    wire N__36646;
    wire N__36641;
    wire N__36632;
    wire N__36623;
    wire N__36614;
    wire N__36609;
    wire N__36606;
    wire N__36601;
    wire N__36598;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36571;
    wire N__36568;
    wire N__36565;
    wire N__36556;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36541;
    wire N__36538;
    wire N__36535;
    wire N__36534;
    wire N__36531;
    wire N__36528;
    wire N__36525;
    wire N__36520;
    wire N__36517;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36486;
    wire N__36481;
    wire N__36478;
    wire N__36477;
    wire N__36474;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36451;
    wire N__36448;
    wire N__36447;
    wire N__36444;
    wire N__36439;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36424;
    wire N__36421;
    wire N__36420;
    wire N__36419;
    wire N__36414;
    wire N__36411;
    wire N__36408;
    wire N__36403;
    wire N__36400;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36387;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36373;
    wire N__36370;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36355;
    wire N__36352;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36337;
    wire N__36334;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36319;
    wire N__36316;
    wire N__36315;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36292;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36277;
    wire N__36274;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36259;
    wire N__36256;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36229;
    wire N__36228;
    wire N__36225;
    wire N__36224;
    wire N__36223;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36209;
    wire N__36206;
    wire N__36201;
    wire N__36198;
    wire N__36195;
    wire N__36190;
    wire N__36189;
    wire N__36184;
    wire N__36181;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36163;
    wire N__36160;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36142;
    wire N__36141;
    wire N__36140;
    wire N__36137;
    wire N__36132;
    wire N__36129;
    wire N__36126;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36116;
    wire N__36109;
    wire N__36106;
    wire N__36103;
    wire N__36100;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36088;
    wire N__36085;
    wire N__36082;
    wire N__36079;
    wire N__36078;
    wire N__36075;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36049;
    wire N__36048;
    wire N__36045;
    wire N__36042;
    wire N__36039;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36007;
    wire N__36004;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35989;
    wire N__35986;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35971;
    wire N__35968;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35949;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35932;
    wire N__35931;
    wire N__35926;
    wire N__35923;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35913;
    wire N__35908;
    wire N__35905;
    wire N__35904;
    wire N__35901;
    wire N__35898;
    wire N__35895;
    wire N__35890;
    wire N__35887;
    wire N__35884;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35873;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35845;
    wire N__35844;
    wire N__35843;
    wire N__35838;
    wire N__35835;
    wire N__35832;
    wire N__35829;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35784;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35772;
    wire N__35769;
    wire N__35766;
    wire N__35761;
    wire N__35758;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35740;
    wire N__35737;
    wire N__35734;
    wire N__35733;
    wire N__35730;
    wire N__35727;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35715;
    wire N__35714;
    wire N__35711;
    wire N__35708;
    wire N__35707;
    wire N__35704;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35676;
    wire N__35675;
    wire N__35674;
    wire N__35671;
    wire N__35668;
    wire N__35663;
    wire N__35656;
    wire N__35655;
    wire N__35652;
    wire N__35651;
    wire N__35650;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35635;
    wire N__35634;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35617;
    wire N__35608;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35587;
    wire N__35584;
    wire N__35583;
    wire N__35580;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35563;
    wire N__35560;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35548;
    wire N__35545;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35514;
    wire N__35511;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35494;
    wire N__35491;
    wire N__35490;
    wire N__35487;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35470;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35458;
    wire N__35457;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35447;
    wire N__35446;
    wire N__35443;
    wire N__35442;
    wire N__35439;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35422;
    wire N__35419;
    wire N__35414;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35382;
    wire N__35379;
    wire N__35376;
    wire N__35373;
    wire N__35370;
    wire N__35367;
    wire N__35366;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35348;
    wire N__35341;
    wire N__35340;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35307;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35284;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35266;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35256;
    wire N__35251;
    wire N__35248;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35211;
    wire N__35208;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35191;
    wire N__35190;
    wire N__35187;
    wire N__35184;
    wire N__35183;
    wire N__35180;
    wire N__35177;
    wire N__35174;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35159;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35123;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35111;
    wire N__35108;
    wire N__35105;
    wire N__35104;
    wire N__35103;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35080;
    wire N__35079;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35069;
    wire N__35062;
    wire N__35059;
    wire N__35056;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35040;
    wire N__35037;
    wire N__35036;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35020;
    wire N__35019;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34983;
    wire N__34980;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34970;
    wire N__34963;
    wire N__34962;
    wire N__34961;
    wire N__34958;
    wire N__34957;
    wire N__34950;
    wire N__34947;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34935;
    wire N__34934;
    wire N__34931;
    wire N__34926;
    wire N__34921;
    wire N__34920;
    wire N__34919;
    wire N__34918;
    wire N__34915;
    wire N__34910;
    wire N__34907;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34891;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34879;
    wire N__34878;
    wire N__34877;
    wire N__34874;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34852;
    wire N__34851;
    wire N__34850;
    wire N__34849;
    wire N__34844;
    wire N__34841;
    wire N__34838;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34787;
    wire N__34784;
    wire N__34779;
    wire N__34776;
    wire N__34775;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34763;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34746;
    wire N__34743;
    wire N__34740;
    wire N__34735;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34723;
    wire N__34720;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34705;
    wire N__34702;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34684;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34660;
    wire N__34659;
    wire N__34656;
    wire N__34653;
    wire N__34650;
    wire N__34649;
    wire N__34646;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34630;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34609;
    wire N__34608;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34598;
    wire N__34597;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34576;
    wire N__34573;
    wire N__34572;
    wire N__34571;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34551;
    wire N__34546;
    wire N__34543;
    wire N__34540;
    wire N__34537;
    wire N__34534;
    wire N__34533;
    wire N__34532;
    wire N__34529;
    wire N__34524;
    wire N__34519;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34507;
    wire N__34506;
    wire N__34505;
    wire N__34502;
    wire N__34497;
    wire N__34492;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34471;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34459;
    wire N__34456;
    wire N__34455;
    wire N__34454;
    wire N__34451;
    wire N__34446;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34408;
    wire N__34405;
    wire N__34402;
    wire N__34399;
    wire N__34396;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34173;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34158;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34140;
    wire N__34139;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34125;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34110;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34100;
    wire N__34097;
    wire N__34090;
    wire N__34087;
    wire N__34086;
    wire N__34085;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34075;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34061;
    wire N__34060;
    wire N__34057;
    wire N__34052;
    wire N__34049;
    wire N__34042;
    wire N__34039;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34012;
    wire N__34011;
    wire N__34008;
    wire N__34007;
    wire N__34006;
    wire N__34003;
    wire N__34002;
    wire N__33999;
    wire N__33994;
    wire N__33989;
    wire N__33984;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33952;
    wire N__33951;
    wire N__33950;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33937;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33918;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33867;
    wire N__33864;
    wire N__33863;
    wire N__33862;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33840;
    wire N__33837;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33817;
    wire N__33814;
    wire N__33813;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33781;
    wire N__33778;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33743;
    wire N__33740;
    wire N__33737;
    wire N__33734;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33717;
    wire N__33716;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33703;
    wire N__33702;
    wire N__33699;
    wire N__33696;
    wire N__33693;
    wire N__33688;
    wire N__33685;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33546;
    wire N__33545;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33478;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33366;
    wire N__33361;
    wire N__33358;
    wire N__33357;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33347;
    wire N__33342;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33312;
    wire N__33309;
    wire N__33306;
    wire N__33303;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33149;
    wire N__33144;
    wire N__33141;
    wire N__33140;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33128;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33087;
    wire N__33086;
    wire N__33085;
    wire N__33084;
    wire N__33081;
    wire N__33072;
    wire N__33067;
    wire N__33066;
    wire N__33063;
    wire N__33062;
    wire N__33061;
    wire N__33056;
    wire N__33053;
    wire N__33050;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32892;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32881;
    wire N__32878;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32857;
    wire N__32854;
    wire N__32853;
    wire N__32852;
    wire N__32851;
    wire N__32850;
    wire N__32849;
    wire N__32848;
    wire N__32845;
    wire N__32842;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32828;
    wire N__32827;
    wire N__32826;
    wire N__32825;
    wire N__32824;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32790;
    wire N__32787;
    wire N__32778;
    wire N__32775;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32740;
    wire N__32737;
    wire N__32734;
    wire N__32731;
    wire N__32728;
    wire N__32727;
    wire N__32726;
    wire N__32725;
    wire N__32724;
    wire N__32723;
    wire N__32722;
    wire N__32721;
    wire N__32720;
    wire N__32719;
    wire N__32718;
    wire N__32717;
    wire N__32716;
    wire N__32715;
    wire N__32712;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32701;
    wire N__32700;
    wire N__32697;
    wire N__32694;
    wire N__32693;
    wire N__32678;
    wire N__32677;
    wire N__32674;
    wire N__32673;
    wire N__32672;
    wire N__32671;
    wire N__32670;
    wire N__32669;
    wire N__32668;
    wire N__32667;
    wire N__32662;
    wire N__32655;
    wire N__32654;
    wire N__32653;
    wire N__32652;
    wire N__32651;
    wire N__32650;
    wire N__32649;
    wire N__32648;
    wire N__32647;
    wire N__32646;
    wire N__32645;
    wire N__32644;
    wire N__32643;
    wire N__32642;
    wire N__32641;
    wire N__32640;
    wire N__32639;
    wire N__32638;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32622;
    wire N__32619;
    wire N__32610;
    wire N__32607;
    wire N__32606;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32598;
    wire N__32597;
    wire N__32596;
    wire N__32595;
    wire N__32594;
    wire N__32593;
    wire N__32592;
    wire N__32589;
    wire N__32588;
    wire N__32587;
    wire N__32586;
    wire N__32585;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32572;
    wire N__32571;
    wire N__32570;
    wire N__32569;
    wire N__32566;
    wire N__32565;
    wire N__32562;
    wire N__32561;
    wire N__32558;
    wire N__32557;
    wire N__32554;
    wire N__32553;
    wire N__32550;
    wire N__32549;
    wire N__32546;
    wire N__32545;
    wire N__32542;
    wire N__32541;
    wire N__32538;
    wire N__32537;
    wire N__32536;
    wire N__32535;
    wire N__32534;
    wire N__32533;
    wire N__32532;
    wire N__32531;
    wire N__32530;
    wire N__32529;
    wire N__32528;
    wire N__32527;
    wire N__32526;
    wire N__32525;
    wire N__32524;
    wire N__32523;
    wire N__32522;
    wire N__32507;
    wire N__32494;
    wire N__32487;
    wire N__32474;
    wire N__32461;
    wire N__32458;
    wire N__32457;
    wire N__32456;
    wire N__32455;
    wire N__32454;
    wire N__32453;
    wire N__32452;
    wire N__32451;
    wire N__32448;
    wire N__32447;
    wire N__32446;
    wire N__32445;
    wire N__32444;
    wire N__32443;
    wire N__32440;
    wire N__32439;
    wire N__32436;
    wire N__32435;
    wire N__32432;
    wire N__32431;
    wire N__32428;
    wire N__32423;
    wire N__32410;
    wire N__32395;
    wire N__32378;
    wire N__32375;
    wire N__32374;
    wire N__32371;
    wire N__32370;
    wire N__32367;
    wire N__32366;
    wire N__32363;
    wire N__32362;
    wire N__32359;
    wire N__32358;
    wire N__32355;
    wire N__32354;
    wire N__32351;
    wire N__32350;
    wire N__32347;
    wire N__32346;
    wire N__32343;
    wire N__32342;
    wire N__32339;
    wire N__32338;
    wire N__32335;
    wire N__32334;
    wire N__32331;
    wire N__32330;
    wire N__32327;
    wire N__32326;
    wire N__32323;
    wire N__32322;
    wire N__32319;
    wire N__32318;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32288;
    wire N__32281;
    wire N__32278;
    wire N__32261;
    wire N__32250;
    wire N__32233;
    wire N__32216;
    wire N__32199;
    wire N__32186;
    wire N__32183;
    wire N__32158;
    wire N__32157;
    wire N__32156;
    wire N__32155;
    wire N__32148;
    wire N__32147;
    wire N__32146;
    wire N__32143;
    wire N__32142;
    wire N__32141;
    wire N__32140;
    wire N__32139;
    wire N__32138;
    wire N__32137;
    wire N__32136;
    wire N__32135;
    wire N__32134;
    wire N__32133;
    wire N__32132;
    wire N__32129;
    wire N__32128;
    wire N__32125;
    wire N__32124;
    wire N__32123;
    wire N__32122;
    wire N__32121;
    wire N__32120;
    wire N__32119;
    wire N__32118;
    wire N__32117;
    wire N__32116;
    wire N__32115;
    wire N__32114;
    wire N__32113;
    wire N__32112;
    wire N__32111;
    wire N__32110;
    wire N__32109;
    wire N__32108;
    wire N__32107;
    wire N__32096;
    wire N__32093;
    wire N__32092;
    wire N__32091;
    wire N__32090;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32086;
    wire N__32083;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32050;
    wire N__32037;
    wire N__32026;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32018;
    wire N__32017;
    wire N__32016;
    wire N__32015;
    wire N__32014;
    wire N__32011;
    wire N__31994;
    wire N__31993;
    wire N__31992;
    wire N__31991;
    wire N__31990;
    wire N__31989;
    wire N__31988;
    wire N__31987;
    wire N__31986;
    wire N__31985;
    wire N__31982;
    wire N__31977;
    wire N__31968;
    wire N__31965;
    wire N__31964;
    wire N__31963;
    wire N__31962;
    wire N__31961;
    wire N__31960;
    wire N__31959;
    wire N__31958;
    wire N__31957;
    wire N__31956;
    wire N__31953;
    wire N__31952;
    wire N__31951;
    wire N__31950;
    wire N__31949;
    wire N__31946;
    wire N__31933;
    wire N__31928;
    wire N__31913;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31897;
    wire N__31882;
    wire N__31879;
    wire N__31866;
    wire N__31859;
    wire N__31854;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31830;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31804;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31789;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31781;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31767;
    wire N__31764;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31675;
    wire N__31672;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31653;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31619;
    wire N__31612;
    wire N__31609;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31595;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31544;
    wire N__31543;
    wire N__31540;
    wire N__31537;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31521;
    wire N__31516;
    wire N__31513;
    wire N__31512;
    wire N__31509;
    wire N__31508;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31428;
    wire N__31423;
    wire N__31420;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31396;
    wire N__31393;
    wire N__31388;
    wire N__31385;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31352;
    wire N__31351;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31312;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31289;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31267;
    wire N__31266;
    wire N__31263;
    wire N__31262;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31243;
    wire N__31240;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31232;
    wire N__31229;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31211;
    wire N__31208;
    wire N__31203;
    wire N__31198;
    wire N__31195;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31169;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31156;
    wire N__31153;
    wire N__31150;
    wire N__31145;
    wire N__31138;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31130;
    wire N__31127;
    wire N__31124;
    wire N__31121;
    wire N__31116;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31063;
    wire N__31060;
    wire N__31059;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31048;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31029;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30985;
    wire N__30982;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30970;
    wire N__30967;
    wire N__30964;
    wire N__30963;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30923;
    wire N__30920;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30902;
    wire N__30897;
    wire N__30892;
    wire N__30889;
    wire N__30888;
    wire N__30885;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30830;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30809;
    wire N__30806;
    wire N__30799;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30777;
    wire N__30772;
    wire N__30769;
    wire N__30766;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30749;
    wire N__30746;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30736;
    wire N__30733;
    wire N__30728;
    wire N__30723;
    wire N__30718;
    wire N__30715;
    wire N__30714;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30681;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30669;
    wire N__30668;
    wire N__30661;
    wire N__30658;
    wire N__30657;
    wire N__30656;
    wire N__30655;
    wire N__30654;
    wire N__30653;
    wire N__30652;
    wire N__30649;
    wire N__30648;
    wire N__30647;
    wire N__30646;
    wire N__30645;
    wire N__30644;
    wire N__30643;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30631;
    wire N__30630;
    wire N__30625;
    wire N__30624;
    wire N__30623;
    wire N__30622;
    wire N__30621;
    wire N__30620;
    wire N__30619;
    wire N__30618;
    wire N__30617;
    wire N__30616;
    wire N__30615;
    wire N__30612;
    wire N__30597;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30578;
    wire N__30573;
    wire N__30570;
    wire N__30559;
    wire N__30552;
    wire N__30535;
    wire N__30532;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30514;
    wire N__30513;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30495;
    wire N__30490;
    wire N__30487;
    wire N__30486;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30312;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30291;
    wire N__30288;
    wire N__30281;
    wire N__30278;
    wire N__30273;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30261;
    wire N__30258;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30147;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30129;
    wire N__30124;
    wire N__30121;
    wire N__30120;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30094;
    wire N__30091;
    wire N__30090;
    wire N__30087;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30069;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30057;
    wire N__30056;
    wire N__30053;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30037;
    wire N__30034;
    wire N__30033;
    wire N__30032;
    wire N__30029;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30003;
    wire N__30000;
    wire N__29999;
    wire N__29998;
    wire N__29997;
    wire N__29994;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29963;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29916;
    wire N__29913;
    wire N__29912;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29895;
    wire N__29890;
    wire N__29887;
    wire N__29886;
    wire N__29883;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29865;
    wire N__29860;
    wire N__29857;
    wire N__29856;
    wire N__29853;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29843;
    wire N__29842;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29812;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29793;
    wire N__29790;
    wire N__29789;
    wire N__29786;
    wire N__29785;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29770;
    wire N__29767;
    wire N__29760;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29718;
    wire N__29715;
    wire N__29714;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29704;
    wire N__29703;
    wire N__29700;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29682;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29641;
    wire N__29638;
    wire N__29637;
    wire N__29634;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29623;
    wire N__29620;
    wire N__29615;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29583;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29483;
    wire N__29482;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29455;
    wire N__29452;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29420;
    wire N__29417;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29373;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29361;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29339;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29297;
    wire N__29290;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29262;
    wire N__29261;
    wire N__29258;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29234;
    wire N__29229;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29204;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29193;
    wire N__29190;
    wire N__29183;
    wire N__29180;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29158;
    wire N__29155;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29143;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29115;
    wire N__29114;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29096;
    wire N__29089;
    wire N__29088;
    wire N__29087;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29048;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29020;
    wire N__29019;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28998;
    wire N__28997;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28938;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28920;
    wire N__28919;
    wire N__28918;
    wire N__28909;
    wire N__28906;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28882;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28870;
    wire N__28869;
    wire N__28866;
    wire N__28863;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28848;
    wire N__28845;
    wire N__28842;
    wire N__28837;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28815;
    wire N__28812;
    wire N__28809;
    wire N__28804;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28771;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28731;
    wire N__28726;
    wire N__28723;
    wire N__28720;
    wire N__28719;
    wire N__28718;
    wire N__28715;
    wire N__28712;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28696;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28662;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28647;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28438;
    wire N__28435;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28410;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28314;
    wire N__28313;
    wire N__28312;
    wire N__28311;
    wire N__28310;
    wire N__28309;
    wire N__28308;
    wire N__28305;
    wire N__28304;
    wire N__28303;
    wire N__28302;
    wire N__28301;
    wire N__28300;
    wire N__28297;
    wire N__28290;
    wire N__28289;
    wire N__28288;
    wire N__28287;
    wire N__28286;
    wire N__28285;
    wire N__28284;
    wire N__28283;
    wire N__28282;
    wire N__28281;
    wire N__28278;
    wire N__28277;
    wire N__28276;
    wire N__28275;
    wire N__28274;
    wire N__28273;
    wire N__28272;
    wire N__28271;
    wire N__28270;
    wire N__28269;
    wire N__28268;
    wire N__28267;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28245;
    wire N__28240;
    wire N__28237;
    wire N__28230;
    wire N__28221;
    wire N__28220;
    wire N__28213;
    wire N__28212;
    wire N__28211;
    wire N__28208;
    wire N__28207;
    wire N__28204;
    wire N__28203;
    wire N__28200;
    wire N__28199;
    wire N__28196;
    wire N__28195;
    wire N__28192;
    wire N__28191;
    wire N__28188;
    wire N__28187;
    wire N__28184;
    wire N__28183;
    wire N__28180;
    wire N__28179;
    wire N__28176;
    wire N__28175;
    wire N__28172;
    wire N__28171;
    wire N__28168;
    wire N__28167;
    wire N__28166;
    wire N__28165;
    wire N__28164;
    wire N__28161;
    wire N__28158;
    wire N__28153;
    wire N__28150;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28132;
    wire N__28117;
    wire N__28100;
    wire N__28083;
    wire N__28082;
    wire N__28079;
    wire N__28078;
    wire N__28075;
    wire N__28074;
    wire N__28071;
    wire N__28070;
    wire N__28067;
    wire N__28062;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28041;
    wire N__28026;
    wire N__28019;
    wire N__28016;
    wire N__28007;
    wire N__28000;
    wire N__27997;
    wire N__27996;
    wire N__27995;
    wire N__27992;
    wire N__27991;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27976;
    wire N__27973;
    wire N__27972;
    wire N__27969;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27943;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27925;
    wire N__27924;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27912;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27882;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27676;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27659;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27634;
    wire N__27633;
    wire N__27632;
    wire N__27631;
    wire N__27630;
    wire N__27629;
    wire N__27628;
    wire N__27627;
    wire N__27626;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27600;
    wire N__27599;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27574;
    wire N__27571;
    wire N__27570;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27558;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27548;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27528;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27518;
    wire N__27515;
    wire N__27512;
    wire N__27509;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27492;
    wire N__27487;
    wire N__27486;
    wire N__27485;
    wire N__27482;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27422;
    wire N__27419;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27401;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27335;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27314;
    wire N__27311;
    wire N__27304;
    wire N__27303;
    wire N__27300;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27280;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27268;
    wire N__27267;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27238;
    wire N__27235;
    wire N__27234;
    wire N__27229;
    wire N__27226;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27189;
    wire N__27186;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27175;
    wire N__27172;
    wire N__27167;
    wire N__27164;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27133;
    wire N__27130;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27093;
    wire N__27092;
    wire N__27089;
    wire N__27084;
    wire N__27079;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27034;
    wire N__27031;
    wire N__27028;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26881;
    wire N__26878;
    wire N__26875;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26541;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26481;
    wire N__26478;
    wire N__26475;
    wire N__26474;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26456;
    wire N__26451;
    wire N__26446;
    wire N__26443;
    wire N__26442;
    wire N__26439;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26419;
    wire N__26416;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26376;
    wire N__26373;
    wire N__26370;
    wire N__26369;
    wire N__26368;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26349;
    wire N__26346;
    wire N__26341;
    wire N__26338;
    wire N__26337;
    wire N__26334;
    wire N__26331;
    wire N__26330;
    wire N__26325;
    wire N__26322;
    wire N__26319;
    wire N__26314;
    wire N__26311;
    wire N__26310;
    wire N__26307;
    wire N__26304;
    wire N__26303;
    wire N__26302;
    wire N__26299;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26282;
    wire N__26279;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26265;
    wire N__26262;
    wire N__26259;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26244;
    wire N__26241;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26223;
    wire N__26220;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26207;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26195;
    wire N__26190;
    wire N__26185;
    wire N__26182;
    wire N__26181;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26140;
    wire N__26137;
    wire N__26134;
    wire N__26133;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26123;
    wire N__26118;
    wire N__26113;
    wire N__26112;
    wire N__26109;
    wire N__26106;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26094;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26077;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26066;
    wire N__26065;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26037;
    wire N__26032;
    wire N__26029;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__25999;
    wire N__25996;
    wire N__25995;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25980;
    wire N__25975;
    wire N__25972;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25958;
    wire N__25953;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25940;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25924;
    wire N__25923;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25879;
    wire N__25876;
    wire N__25875;
    wire N__25872;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25827;
    wire N__25826;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25808;
    wire N__25803;
    wire N__25798;
    wire N__25795;
    wire N__25794;
    wire N__25791;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25557;
    wire N__25556;
    wire N__25555;
    wire N__25554;
    wire N__25553;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25547;
    wire N__25546;
    wire N__25543;
    wire N__25542;
    wire N__25539;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25531;
    wire N__25528;
    wire N__25527;
    wire N__25524;
    wire N__25523;
    wire N__25520;
    wire N__25519;
    wire N__25518;
    wire N__25501;
    wire N__25484;
    wire N__25481;
    wire N__25480;
    wire N__25475;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25390;
    wire N__25387;
    wire N__25384;
    wire N__25381;
    wire N__25380;
    wire N__25379;
    wire N__25376;
    wire N__25375;
    wire N__25372;
    wire N__25369;
    wire N__25366;
    wire N__25363;
    wire N__25360;
    wire N__25357;
    wire N__25350;
    wire N__25345;
    wire N__25344;
    wire N__25343;
    wire N__25342;
    wire N__25333;
    wire N__25332;
    wire N__25331;
    wire N__25330;
    wire N__25329;
    wire N__25328;
    wire N__25327;
    wire N__25326;
    wire N__25325;
    wire N__25324;
    wire N__25323;
    wire N__25322;
    wire N__25321;
    wire N__25320;
    wire N__25319;
    wire N__25318;
    wire N__25317;
    wire N__25316;
    wire N__25315;
    wire N__25314;
    wire N__25313;
    wire N__25312;
    wire N__25311;
    wire N__25310;
    wire N__25309;
    wire N__25308;
    wire N__25307;
    wire N__25304;
    wire N__25295;
    wire N__25286;
    wire N__25277;
    wire N__25272;
    wire N__25263;
    wire N__25254;
    wire N__25245;
    wire N__25240;
    wire N__25235;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24954;
    wire N__24953;
    wire N__24946;
    wire N__24943;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24925;
    wire N__24922;
    wire N__24921;
    wire N__24916;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24904;
    wire N__24901;
    wire N__24900;
    wire N__24899;
    wire N__24896;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24859;
    wire N__24858;
    wire N__24855;
    wire N__24854;
    wire N__24851;
    wire N__24848;
    wire N__24845;
    wire N__24838;
    wire N__24835;
    wire N__24834;
    wire N__24833;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24817;
    wire N__24814;
    wire N__24813;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24802;
    wire N__24795;
    wire N__24792;
    wire N__24787;
    wire N__24786;
    wire N__24783;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24771;
    wire N__24768;
    wire N__24763;
    wire N__24762;
    wire N__24757;
    wire N__24756;
    wire N__24753;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24724;
    wire N__24723;
    wire N__24720;
    wire N__24715;
    wire N__24712;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24688;
    wire N__24687;
    wire N__24684;
    wire N__24683;
    wire N__24680;
    wire N__24675;
    wire N__24672;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24570;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24553;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24504;
    wire N__24503;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24489;
    wire N__24484;
    wire N__24481;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24459;
    wire N__24454;
    wire N__24451;
    wire N__24450;
    wire N__24449;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24426;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24411;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24351;
    wire N__24350;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24334;
    wire N__24331;
    wire N__24328;
    wire N__24327;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24312;
    wire N__24307;
    wire N__24304;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24282;
    wire N__24277;
    wire N__24274;
    wire N__24273;
    wire N__24272;
    wire N__24267;
    wire N__24264;
    wire N__24261;
    wire N__24256;
    wire N__24253;
    wire N__24250;
    wire N__24249;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24234;
    wire N__24229;
    wire N__24226;
    wire N__24225;
    wire N__24222;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24207;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24195;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24180;
    wire N__24175;
    wire N__24172;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24164;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24148;
    wire N__24145;
    wire N__24144;
    wire N__24143;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24127;
    wire N__24124;
    wire N__24123;
    wire N__24122;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24106;
    wire N__24103;
    wire N__24100;
    wire N__24099;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24084;
    wire N__24079;
    wire N__24076;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24051;
    wire N__24046;
    wire N__24043;
    wire N__24042;
    wire N__24041;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24018;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24003;
    wire N__23998;
    wire N__23995;
    wire N__23994;
    wire N__23991;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23976;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23964;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23949;
    wire N__23944;
    wire N__23941;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23933;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23917;
    wire N__23914;
    wire N__23913;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23886;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23871;
    wire N__23866;
    wire N__23863;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23855;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23839;
    wire N__23836;
    wire N__23835;
    wire N__23832;
    wire N__23829;
    wire N__23828;
    wire N__23823;
    wire N__23820;
    wire N__23817;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23805;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23790;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23778;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23763;
    wire N__23758;
    wire N__23755;
    wire N__23752;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23744;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23689;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23407;
    wire N__23404;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23338;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23278;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23244;
    wire N__23241;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23193;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23175;
    wire N__23172;
    wire N__23171;
    wire N__23170;
    wire N__23169;
    wire N__23168;
    wire N__23167;
    wire N__23166;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23150;
    wire N__23143;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23119;
    wire N__23114;
    wire N__23111;
    wire N__23108;
    wire N__23105;
    wire N__23098;
    wire N__23095;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23032;
    wire N__23029;
    wire N__23028;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23013;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22995;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22959;
    wire N__22956;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22872;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22828;
    wire N__22825;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22804;
    wire N__22801;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22780;
    wire N__22777;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22729;
    wire N__22726;
    wire N__22725;
    wire N__22724;
    wire N__22721;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22692;
    wire N__22691;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22679;
    wire N__22676;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22623;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22608;
    wire N__22607;
    wire N__22604;
    wire N__22601;
    wire N__22598;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22582;
    wire N__22579;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22551;
    wire N__22546;
    wire N__22543;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22525;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22503;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22479;
    wire N__22474;
    wire N__22471;
    wire N__22470;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22383;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22363;
    wire N__22360;
    wire N__22359;
    wire N__22358;
    wire N__22357;
    wire N__22356;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22335;
    wire N__22330;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22312;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22266;
    wire N__22261;
    wire N__22258;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22223;
    wire N__22218;
    wire N__22215;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22198;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22175;
    wire N__22174;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22156;
    wire N__22153;
    wire N__22148;
    wire N__22145;
    wire N__22138;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22123;
    wire N__22122;
    wire N__22121;
    wire N__22120;
    wire N__22119;
    wire N__22118;
    wire N__22115;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22096;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22081;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22059;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22015;
    wire N__22014;
    wire N__22013;
    wire N__22010;
    wire N__22009;
    wire N__22006;
    wire N__22005;
    wire N__22004;
    wire N__22003;
    wire N__22000;
    wire N__21999;
    wire N__21998;
    wire N__21991;
    wire N__21988;
    wire N__21985;
    wire N__21982;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21968;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21948;
    wire N__21945;
    wire N__21940;
    wire N__21929;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21915;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21880;
    wire N__21879;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21844;
    wire N__21841;
    wire N__21840;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21825;
    wire N__21822;
    wire N__21817;
    wire N__21814;
    wire N__21813;
    wire N__21808;
    wire N__21807;
    wire N__21806;
    wire N__21805;
    wire N__21804;
    wire N__21803;
    wire N__21802;
    wire N__21801;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21779;
    wire N__21774;
    wire N__21769;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21761;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21745;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21723;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21699;
    wire N__21696;
    wire N__21691;
    wire N__21690;
    wire N__21687;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21669;
    wire N__21666;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21648;
    wire N__21645;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21606;
    wire N__21605;
    wire N__21604;
    wire N__21603;
    wire N__21602;
    wire N__21601;
    wire N__21600;
    wire N__21599;
    wire N__21598;
    wire N__21583;
    wire N__21580;
    wire N__21575;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21432;
    wire N__21431;
    wire N__21430;
    wire N__21429;
    wire N__21428;
    wire N__21425;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21419;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21411;
    wire N__21410;
    wire N__21409;
    wire N__21408;
    wire N__21407;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21382;
    wire N__21379;
    wire N__21378;
    wire N__21373;
    wire N__21366;
    wire N__21361;
    wire N__21356;
    wire N__21355;
    wire N__21354;
    wire N__21353;
    wire N__21352;
    wire N__21351;
    wire N__21350;
    wire N__21349;
    wire N__21348;
    wire N__21347;
    wire N__21346;
    wire N__21345;
    wire N__21344;
    wire N__21343;
    wire N__21342;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21330;
    wire N__21325;
    wire N__21308;
    wire N__21293;
    wire N__21286;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21205;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21197;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21181;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21046;
    wire N__21045;
    wire N__21042;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21013;
    wire N__21012;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20997;
    wire N__20992;
    wire N__20989;
    wire N__20986;
    wire N__20985;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20972;
    wire N__20969;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20952;
    wire N__20949;
    wire N__20948;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20932;
    wire N__20929;
    wire N__20926;
    wire N__20925;
    wire N__20922;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20896;
    wire N__20893;
    wire N__20890;
    wire N__20887;
    wire N__20884;
    wire N__20881;
    wire N__20878;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20838;
    wire N__20835;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20820;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20808;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20793;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20762;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20739;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20724;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20700;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20685;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20673;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20658;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20544;
    wire N__20541;
    wire N__20538;
    wire N__20535;
    wire N__20532;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20355;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20331;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20281;
    wire N__20280;
    wire N__20275;
    wire N__20272;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20242;
    wire N__20239;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20217;
    wire N__20216;
    wire N__20213;
    wire N__20208;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20196;
    wire N__20193;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20007;
    wire N__20006;
    wire N__20005;
    wire N__20004;
    wire N__20003;
    wire N__20002;
    wire N__20001;
    wire N__20000;
    wire N__19999;
    wire N__19990;
    wire N__19981;
    wire N__19976;
    wire N__19971;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19846;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19776;
    wire N__19775;
    wire N__19774;
    wire N__19773;
    wire N__19772;
    wire N__19769;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19741;
    wire N__19732;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire bfn_1_11_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire bfn_1_12_0_;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire bfn_1_13_0_;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire N_42_i_i;
    wire un7_start_stop_0_a2;
    wire bfn_2_5_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_2_6_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_2_8_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_2_9_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire bfn_2_10_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10_cascade_ ;
    wire pwm_duty_input_1;
    wire pwm_duty_input_0;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12_cascade_ ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13_cascade_ ;
    wire \pwm_generator_inst.un3_threshold ;
    wire bfn_2_13_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ;
    wire bfn_2_14_0_;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0 ;
    wire bfn_2_15_0_;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_3_7_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_3_8_0_;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire bfn_3_9_0_;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire bfn_3_10_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8 ;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.N_149 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31 ;
    wire \pwm_generator_inst.threshold_0 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671 ;
    wire \pwm_generator_inst.threshold_9 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791 ;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61 ;
    wire N_19_1;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_6;
    wire pwm_duty_input_8;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ;
    wire \pwm_generator_inst.N_17 ;
    wire \current_shift_inst.PI_CTRL.N_154 ;
    wire pwm_duty_input_2;
    wire pwm_duty_input_7;
    wire pwm_duty_input_5;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire pwm_duty_input_4;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \pwm_generator_inst.N_16 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_53_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.N_155 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire delay_hc_input_c_g;
    wire il_max_comp2_c;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ;
    wire \current_shift_inst.PI_CTRL.N_153 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.N_53 ;
    wire pwm_duty_input_3;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire bfn_7_9_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire bfn_7_10_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire bfn_7_11_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire bfn_7_12_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire bfn_7_19_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_7_20_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_7_21_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_7_22_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire il_min_comp2_c;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ;
    wire il_max_comp2_D1;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_72_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire bfn_8_13_0_;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire bfn_8_14_0_;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire bfn_8_15_0_;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire bfn_8_16_0_;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_8_21_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_8_22_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_8_23_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_8_24_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire il_min_comp1_c;
    wire il_max_comp1_c;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.un1_enablelt3_0 ;
    wire \current_shift_inst.PI_CTRL.N_71 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire il_min_comp2_D1;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire bfn_9_17_0_;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_9_18_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire bfn_9_20_0_;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire s3_phy_c;
    wire \current_shift_inst.timer_s1.running_i ;
    wire s4_phy_c;
    wire il_max_comp1_D1;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire bfn_10_13_0_;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ;
    wire bfn_10_14_0_;
    wire \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_10_15_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire bfn_10_16_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_397_i ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire bfn_10_22_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_10_23_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_10_24_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_10_25_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire bfn_11_6_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integrator_i_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_7 ;
    wire bfn_11_7_0_;
    wire \current_shift_inst.PI_CTRL.integrator_i_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire bfn_11_8_0_;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire bfn_11_9_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un13_integrator_cry_30 ;
    wire bfn_11_10_0_;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_26 ;
    wire il_min_comp1_D1;
    wire \current_shift_inst.PI_CTRL.integrator_i_23 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.N_166_i_g ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire bfn_11_15_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ;
    wire bfn_11_16_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ;
    wire bfn_11_17_0_;
    wire \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire bfn_11_18_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_11_20_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_11_21_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire bfn_11_22_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df24 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_399_i ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_i_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_12_9_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire bfn_12_10_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.N_1474_i ;
    wire \current_shift_inst.control_input_18 ;
    wire bfn_12_11_0_;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_12_12_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.control_input_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_ ;
    wire elapsed_time_ns_1_RNIRB3CP1_0_3_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire start_stop_c;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.N_54 ;
    wire \current_shift_inst.timer_s1.N_167_i ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ;
    wire bfn_13_4_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_8 ;
    wire bfn_13_5_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ;
    wire bfn_13_6_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ;
    wire bfn_13_7_0_;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_31 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ;
    wire \pll_inst.red_c_i ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_13_13_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_13_14_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire bfn_13_15_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire elapsed_time_ns_1_RNIPKKEE1_0_8;
    wire elapsed_time_ns_1_RNIOJKEE1_0_7_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_330_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_ ;
    wire elapsed_time_ns_1_RNIRB3CP1_0_3;
    wire elapsed_time_ns_1_RNIJEKEE1_0_2;
    wire \phase_controller_inst1.stoper_hc.N_286 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_328_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ;
    wire elapsed_time_ns_1_RNIP93CP1_0_1;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ;
    wire elapsed_time_ns_1_RNIP93CP1_0_1_cascade_;
    wire \phase_controller_inst1.stoper_hc.N_310 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire state_ns_i_a2_1;
    wire \phase_controller_inst1.tr_time_passed ;
    wire T45_c;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire s1_phy_c;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire T23_c;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_166_i ;
    wire s2_phy_c;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_28_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_16 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_i_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ;
    wire elapsed_time_ns_1_RNIP7HF91_0_10_cascade_;
    wire elapsed_time_ns_1_RNIFJ2591_0_7;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_ ;
    wire elapsed_time_ns_1_RNIGK2591_0_8;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire il_min_comp2_D2;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire \phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_14_15_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_14_16_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_14_17_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_14_18_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df22 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df26 ;
    wire elapsed_time_ns_1_RNIOJKEE1_0_7;
    wire il_max_comp1_D2;
    wire state_3;
    wire T01_c;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0 ;
    wire \current_shift_inst.PI_CTRL.N_74 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_75 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire elapsed_time_ns_1_RNIVEIF91_0_25;
    wire elapsed_time_ns_1_RNIVEIF91_0_25_cascade_;
    wire elapsed_time_ns_1_RNI2IIF91_0_28;
    wire elapsed_time_ns_1_RNI1HIF91_0_27;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ;
    wire elapsed_time_ns_1_RNISBIF91_0_22;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ;
    wire elapsed_time_ns_1_RNI0GIF91_0_26;
    wire elapsed_time_ns_1_RNIP7HF91_0_10;
    wire elapsed_time_ns_1_RNIQ8HF91_0_11;
    wire elapsed_time_ns_1_RNIR9HF91_0_12;
    wire elapsed_time_ns_1_RNISAHF91_0_13;
    wire elapsed_time_ns_1_RNIUCHF91_0_15;
    wire elapsed_time_ns_1_RNIUCHF91_0_15_cascade_;
    wire \phase_controller_inst1.stoper_tr.N_244 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ;
    wire \delay_measurement_inst.delay_tr_timer.N_386_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ;
    wire elapsed_time_ns_1_RNIAE2591_0_2;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_ ;
    wire elapsed_time_ns_1_RNII6NQL1_0_1;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ;
    wire elapsed_time_ns_1_RNII6NQL1_0_1_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ;
    wire elapsed_time_ns_1_RNISCJF91_0_31_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_15_13_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_15_14_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire bfn_15_15_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire elapsed_time_ns_1_RNI4HV8E1_0_30;
    wire elapsed_time_ns_1_RNILGKEE1_0_4;
    wire elapsed_time_ns_1_RNILGKEE1_0_4_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2 ;
    wire elapsed_time_ns_1_RNI4GU8E1_0_21;
    wire elapsed_time_ns_1_RNICOU8E1_0_29;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire bfn_15_17_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire bfn_15_18_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_15_19_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_15_20_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire \delay_measurement_inst.delay_hc_timer.N_397_i_g ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_15_21_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_15_22_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_15_23_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_15_24_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_398_i ;
    wire elapsed_time_ns_1_RNIQ9IF91_0_20;
    wire elapsed_time_ns_1_RNIRAIF91_0_21;
    wire elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_;
    wire elapsed_time_ns_1_RNI3JIF91_0_29;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15 ;
    wire elapsed_time_ns_1_RNITCIF91_0_23;
    wire elapsed_time_ns_1_RNITCIF91_0_23_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ;
    wire elapsed_time_ns_1_RNIUDIF91_0_24;
    wire \delay_measurement_inst.delay_tr_timer.N_379_cascade_ ;
    wire \delay_measurement_inst.delay_tr9_cascade_ ;
    wire elapsed_time_ns_1_RNIRBJF91_0_30;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_358 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ;
    wire \delay_measurement_inst.delay_tr_timer.N_354 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ;
    wire elapsed_time_ns_1_RNIK8NQL1_0_3;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6 ;
    wire elapsed_time_ns_1_RNINBNQL1_0_6;
    wire \delay_measurement_inst.delay_tr_timer.N_353 ;
    wire \delay_measurement_inst.delay_tr_timer.N_353_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_382 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ;
    wire elapsed_time_ns_1_RNIDH2591_0_5;
    wire elapsed_time_ns_1_RNIA965M1_0_18_cascade_;
    wire elapsed_time_ns_1_RNICG2591_0_4;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ;
    wire elapsed_time_ns_1_RNI9865M1_0_17_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lt31_0_2 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14 ;
    wire elapsed_time_ns_1_RNI6565M1_0_14;
    wire \delay_measurement_inst.delay_tr_timer.N_395 ;
    wire \delay_measurement_inst.delay_tr_timer.N_375 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ;
    wire elapsed_time_ns_1_RNIQENQL1_0_9;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_ ;
    wire \phase_controller_inst2.state_RNIG7JFZ0Z_2 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire il_max_comp2_D2;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire elapsed_time_ns_1_RNI8765M1_0_16;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire elapsed_time_ns_1_RNI9865M1_0_17;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire elapsed_time_ns_1_RNIBA65M1_0_19;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire elapsed_time_ns_1_RNISCJF91_0_31;
    wire \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ;
    wire elapsed_time_ns_1_RNIA965M1_0_18;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_ ;
    wire elapsed_time_ns_1_RNI4FT8E1_0_12_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_369_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_367_clk_cascade_ ;
    wire elapsed_time_ns_1_RNI3FU8E1_0_20;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire elapsed_time_ns_1_RNIMHKEE1_0_5;
    wire \phase_controller_inst1.stoper_hc.N_330 ;
    wire elapsed_time_ns_1_RNIMHKEE1_0_5_cascade_;
    wire \phase_controller_inst1.stoper_hc.N_328 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire elapsed_time_ns_1_RNIAMU8E1_0_27;
    wire elapsed_time_ns_1_RNI9LU8E1_0_26;
    wire elapsed_time_ns_1_RNIBNU8E1_0_28;
    wire elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_;
    wire elapsed_time_ns_1_RNI8KU8E1_0_25;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15 ;
    wire elapsed_time_ns_1_RNI5HU8E1_0_22;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15_cascade_ ;
    wire elapsed_time_ns_1_RNI7JU8E1_0_24;
    wire elapsed_time_ns_1_RNI6IU8E1_0_23;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire \delay_measurement_inst.delay_hc_timer.N_369 ;
    wire \delay_measurement_inst.delay_hc_timer.N_344_i_cascade_ ;
    wire elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ;
    wire elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_ ;
    wire elapsed_time_ns_1_RNIGGC6P1_0_17;
    wire elapsed_time_ns_1_RNIGGC6P1_0_17_cascade_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire elapsed_time_ns_1_RNIFFC6P1_0_16;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire elapsed_time_ns_1_RNIIIC6P1_0_19;
    wire \phase_controller_inst1.stoper_hc.N_318_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire elapsed_time_ns_1_RNIHHC6P1_0_18;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire elapsed_time_ns_1_RNI2DT8E1_0_10;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire elapsed_time_ns_1_RNI3ET8E1_0_11;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire elapsed_time_ns_1_RNI4FT8E1_0_12;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire bfn_17_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_17_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_17_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_400_i ;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire bfn_17_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_17_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire bfn_17_14_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.elapsed_time_tr_31 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire il_min_comp1_D2;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst1.N_55 ;
    wire \phase_controller_inst1.start_timer_tr_RNOZ0Z_0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire elapsed_time_ns_1_RNI5GT8E1_0_13;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.N_344_i ;
    wire elapsed_time_ns_1_RNIUE3CP1_0_6;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire elapsed_time_ns_1_RNI7IT8E1_0_15_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.N_269_iZ0Z_1 ;
    wire elapsed_time_ns_1_RNI7IT8E1_0_15;
    wire \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire elapsed_time_ns_1_RNI1I3CP1_0_9;
    wire \delay_measurement_inst.delay_hc_timer.N_367_clk ;
    wire \delay_measurement_inst.delay_tr9 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_17_19_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_17_20_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire bfn_17_21_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire elapsed_time_ns_1_RNI5IV8E1_0_31;
    wire \phase_controller_inst1.stoper_hc.N_318 ;
    wire elapsed_time_ns_1_RNIDDC6P1_0_14;
    wire \phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire T12_c;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.N_399_i_g ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_394 ;
    wire \delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.N_346 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire \delay_measurement_inst.delay_tr_timer.N_346_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.N_349 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.N_349_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.N_351 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \delay_measurement_inst.delay_tr_timer.N_362 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ;
    wire \delay_measurement_inst.delay_tr_timer.N_362_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ;
    wire \delay_measurement_inst.N_365 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_18_13_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_18_14_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_18_15_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire bfn_18_16_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire bfn_18_17_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_18_18_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_18_19_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire bfn_18_20_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df22 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df20 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire red_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__21169),
            .RESETB(N__34198),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__28314),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__28300),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({dangling_wire_16,N__21354,N__21347,N__21352,N__21346,N__21353,N__21345,N__21355,N__21342,N__21348,N__21341,N__21349,N__21343,N__21350,N__21344,N__21351}),
            .C({dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32}),
            .B({dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,N__28313,N__28303,dangling_wire_40,dangling_wire_41,dangling_wire_42,N__28301,N__28312,N__28302,N__28311}),
            .OHOLDTOP(),
            .O({dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__28289),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__28282),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73}),
            .ADDSUBBOT(),
            .A({dangling_wire_74,N__21406,N__21409,N__21407,N__21410,N__21408,N__21914,N__21839,N__21722,N__21878,N__21690,N__21644,N__22390,N__21745,N__20257,N__20242}),
            .C({dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90}),
            .B({dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,N__28288,N__28285,dangling_wire_98,dangling_wire_99,dangling_wire_100,N__28283,N__28287,N__28284,N__28286}),
            .OHOLDTOP(),
            .O({dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__50555),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__50557),
            .DIN(N__50556),
            .DOUT(N__50555),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__50557),
            .PADOUT(N__50556),
            .PADIN(N__50555),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__50546),
            .DIN(N__50545),
            .DOUT(N__50544),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__50546),
            .PADOUT(N__50545),
            .PADIN(N__50544),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__38215),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__50537),
            .DIN(N__50536),
            .DOUT(N__50535),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__50537),
            .PADOUT(N__50536),
            .PADIN(N__50535),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__50528),
            .DIN(N__50527),
            .DOUT(N__50526),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__50528),
            .PADOUT(N__50527),
            .PADIN(N__50526),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__50519),
            .DIN(N__50518),
            .DOUT(N__50517),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__50519),
            .PADOUT(N__50518),
            .PADIN(N__50517),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34900),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__50510),
            .DIN(N__50509),
            .DOUT(N__50508),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__50510),
            .PADOUT(N__50509),
            .PADIN(N__50508),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20896),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__50501),
            .DIN(N__50500),
            .DOUT(N__50499),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__50501),
            .PADOUT(N__50500),
            .PADIN(N__50499),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__50492),
            .DIN(N__50491),
            .DOUT(N__50490),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__50492),
            .PADOUT(N__50491),
            .PADIN(N__50490),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34822),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__50483),
            .DIN(N__50482),
            .DOUT(N__50481),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__50483),
            .PADOUT(N__50482),
            .PADIN(N__50481),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__46555),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__50474),
            .DIN(N__50473),
            .DOUT(N__50472),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__50474),
            .PADOUT(N__50473),
            .PADIN(N__50472),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__50465),
            .DIN(N__50464),
            .DOUT(N__50463),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__50465),
            .PADOUT(N__50464),
            .PADIN(N__50463),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34942),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__50456),
            .DIN(N__50455),
            .DOUT(N__50454),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__50456),
            .PADOUT(N__50455),
            .PADIN(N__50454),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25222),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__50447),
            .DIN(N__50446),
            .DOUT(N__50445),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__50447),
            .PADOUT(N__50446),
            .PADIN(N__50445),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__50438),
            .DIN(N__50437),
            .DOUT(N__50436),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__50438),
            .PADOUT(N__50437),
            .PADIN(N__50436),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25132),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__50429),
            .DIN(N__50428),
            .DOUT(N__50427),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__50429),
            .PADOUT(N__50428),
            .PADIN(N__50427),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34630),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__50420),
            .DIN(N__50419),
            .DOUT(N__50418),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__50420),
            .PADOUT(N__50419),
            .PADIN(N__50418),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__50411),
            .DIN(N__50410),
            .DOUT(N__50409),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__50411),
            .PADOUT(N__50410),
            .PADIN(N__50409),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11955 (
            .O(N__50392),
            .I(N__50388));
    InMux I__11954 (
            .O(N__50391),
            .I(N__50385));
    LocalMux I__11953 (
            .O(N__50388),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__11952 (
            .O(N__50385),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__11951 (
            .O(N__50380),
            .I(N__50376));
    InMux I__11950 (
            .O(N__50379),
            .I(N__50373));
    LocalMux I__11949 (
            .O(N__50376),
            .I(N__50370));
    LocalMux I__11948 (
            .O(N__50373),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__11947 (
            .O(N__50370),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__11946 (
            .O(N__50365),
            .I(N__50362));
    LocalMux I__11945 (
            .O(N__50362),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df24 ));
    InMux I__11944 (
            .O(N__50359),
            .I(N__50355));
    InMux I__11943 (
            .O(N__50358),
            .I(N__50352));
    LocalMux I__11942 (
            .O(N__50355),
            .I(N__50349));
    LocalMux I__11941 (
            .O(N__50352),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__11940 (
            .O(N__50349),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__11939 (
            .O(N__50344),
            .I(N__50340));
    InMux I__11938 (
            .O(N__50343),
            .I(N__50337));
    LocalMux I__11937 (
            .O(N__50340),
            .I(N__50334));
    LocalMux I__11936 (
            .O(N__50337),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__11935 (
            .O(N__50334),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__11934 (
            .O(N__50329),
            .I(N__50326));
    LocalMux I__11933 (
            .O(N__50326),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df20 ));
    CEMux I__11932 (
            .O(N__50323),
            .I(N__50317));
    CEMux I__11931 (
            .O(N__50322),
            .I(N__50314));
    CEMux I__11930 (
            .O(N__50321),
            .I(N__50311));
    CEMux I__11929 (
            .O(N__50320),
            .I(N__50308));
    LocalMux I__11928 (
            .O(N__50317),
            .I(N__50296));
    LocalMux I__11927 (
            .O(N__50314),
            .I(N__50296));
    LocalMux I__11926 (
            .O(N__50311),
            .I(N__50285));
    LocalMux I__11925 (
            .O(N__50308),
            .I(N__50266));
    InMux I__11924 (
            .O(N__50307),
            .I(N__50259));
    InMux I__11923 (
            .O(N__50306),
            .I(N__50259));
    InMux I__11922 (
            .O(N__50305),
            .I(N__50259));
    InMux I__11921 (
            .O(N__50304),
            .I(N__50250));
    InMux I__11920 (
            .O(N__50303),
            .I(N__50250));
    InMux I__11919 (
            .O(N__50302),
            .I(N__50250));
    InMux I__11918 (
            .O(N__50301),
            .I(N__50250));
    Span4Mux_v I__11917 (
            .O(N__50296),
            .I(N__50247));
    InMux I__11916 (
            .O(N__50295),
            .I(N__50240));
    InMux I__11915 (
            .O(N__50294),
            .I(N__50240));
    InMux I__11914 (
            .O(N__50293),
            .I(N__50240));
    InMux I__11913 (
            .O(N__50292),
            .I(N__50237));
    InMux I__11912 (
            .O(N__50291),
            .I(N__50228));
    InMux I__11911 (
            .O(N__50290),
            .I(N__50228));
    InMux I__11910 (
            .O(N__50289),
            .I(N__50228));
    InMux I__11909 (
            .O(N__50288),
            .I(N__50228));
    Span4Mux_v I__11908 (
            .O(N__50285),
            .I(N__50225));
    InMux I__11907 (
            .O(N__50284),
            .I(N__50216));
    InMux I__11906 (
            .O(N__50283),
            .I(N__50216));
    InMux I__11905 (
            .O(N__50282),
            .I(N__50216));
    InMux I__11904 (
            .O(N__50281),
            .I(N__50216));
    InMux I__11903 (
            .O(N__50280),
            .I(N__50207));
    InMux I__11902 (
            .O(N__50279),
            .I(N__50207));
    InMux I__11901 (
            .O(N__50278),
            .I(N__50207));
    InMux I__11900 (
            .O(N__50277),
            .I(N__50207));
    InMux I__11899 (
            .O(N__50276),
            .I(N__50198));
    InMux I__11898 (
            .O(N__50275),
            .I(N__50198));
    InMux I__11897 (
            .O(N__50274),
            .I(N__50198));
    InMux I__11896 (
            .O(N__50273),
            .I(N__50198));
    InMux I__11895 (
            .O(N__50272),
            .I(N__50189));
    InMux I__11894 (
            .O(N__50271),
            .I(N__50189));
    InMux I__11893 (
            .O(N__50270),
            .I(N__50189));
    InMux I__11892 (
            .O(N__50269),
            .I(N__50189));
    Span4Mux_v I__11891 (
            .O(N__50266),
            .I(N__50184));
    LocalMux I__11890 (
            .O(N__50259),
            .I(N__50184));
    LocalMux I__11889 (
            .O(N__50250),
            .I(N__50181));
    Span4Mux_h I__11888 (
            .O(N__50247),
            .I(N__50172));
    LocalMux I__11887 (
            .O(N__50240),
            .I(N__50172));
    LocalMux I__11886 (
            .O(N__50237),
            .I(N__50172));
    LocalMux I__11885 (
            .O(N__50228),
            .I(N__50172));
    Span4Mux_h I__11884 (
            .O(N__50225),
            .I(N__50165));
    LocalMux I__11883 (
            .O(N__50216),
            .I(N__50165));
    LocalMux I__11882 (
            .O(N__50207),
            .I(N__50165));
    LocalMux I__11881 (
            .O(N__50198),
            .I(N__50160));
    LocalMux I__11880 (
            .O(N__50189),
            .I(N__50160));
    Span4Mux_h I__11879 (
            .O(N__50184),
            .I(N__50155));
    Span4Mux_h I__11878 (
            .O(N__50181),
            .I(N__50155));
    Span4Mux_h I__11877 (
            .O(N__50172),
            .I(N__50152));
    Span4Mux_h I__11876 (
            .O(N__50165),
            .I(N__50149));
    Odrv4 I__11875 (
            .O(N__50160),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11874 (
            .O(N__50155),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11873 (
            .O(N__50152),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11872 (
            .O(N__50149),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__11871 (
            .O(N__50140),
            .I(N__50136));
    InMux I__11870 (
            .O(N__50139),
            .I(N__50133));
    LocalMux I__11869 (
            .O(N__50136),
            .I(N__50128));
    LocalMux I__11868 (
            .O(N__50133),
            .I(N__50125));
    InMux I__11867 (
            .O(N__50132),
            .I(N__50122));
    InMux I__11866 (
            .O(N__50131),
            .I(N__50119));
    Span4Mux_v I__11865 (
            .O(N__50128),
            .I(N__50112));
    Span4Mux_v I__11864 (
            .O(N__50125),
            .I(N__50112));
    LocalMux I__11863 (
            .O(N__50122),
            .I(N__50112));
    LocalMux I__11862 (
            .O(N__50119),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__11861 (
            .O(N__50112),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__11860 (
            .O(N__50107),
            .I(N__50103));
    InMux I__11859 (
            .O(N__50106),
            .I(N__50099));
    LocalMux I__11858 (
            .O(N__50103),
            .I(N__50095));
    InMux I__11857 (
            .O(N__50102),
            .I(N__50092));
    LocalMux I__11856 (
            .O(N__50099),
            .I(N__50089));
    InMux I__11855 (
            .O(N__50098),
            .I(N__50085));
    Span12Mux_h I__11854 (
            .O(N__50095),
            .I(N__50082));
    LocalMux I__11853 (
            .O(N__50092),
            .I(N__50079));
    Span4Mux_v I__11852 (
            .O(N__50089),
            .I(N__50076));
    InMux I__11851 (
            .O(N__50088),
            .I(N__50073));
    LocalMux I__11850 (
            .O(N__50085),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv12 I__11849 (
            .O(N__50082),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__11848 (
            .O(N__50079),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__11847 (
            .O(N__50076),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__11846 (
            .O(N__50073),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__11845 (
            .O(N__50062),
            .I(N__50059));
    LocalMux I__11844 (
            .O(N__50059),
            .I(N__50055));
    InMux I__11843 (
            .O(N__50058),
            .I(N__50052));
    Span4Mux_h I__11842 (
            .O(N__50055),
            .I(N__50049));
    LocalMux I__11841 (
            .O(N__50052),
            .I(N__50046));
    Span4Mux_h I__11840 (
            .O(N__50049),
            .I(N__50041));
    Span4Mux_h I__11839 (
            .O(N__50046),
            .I(N__50041));
    Odrv4 I__11838 (
            .O(N__50041),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    CascadeMux I__11837 (
            .O(N__50038),
            .I(N__50034));
    CascadeMux I__11836 (
            .O(N__50037),
            .I(N__50031));
    InMux I__11835 (
            .O(N__50034),
            .I(N__50028));
    InMux I__11834 (
            .O(N__50031),
            .I(N__50025));
    LocalMux I__11833 (
            .O(N__50028),
            .I(N__50022));
    LocalMux I__11832 (
            .O(N__50025),
            .I(N__50019));
    Span4Mux_v I__11831 (
            .O(N__50022),
            .I(N__50011));
    Span4Mux_v I__11830 (
            .O(N__50019),
            .I(N__50011));
    InMux I__11829 (
            .O(N__50018),
            .I(N__50006));
    InMux I__11828 (
            .O(N__50017),
            .I(N__50006));
    InMux I__11827 (
            .O(N__50016),
            .I(N__50003));
    Sp12to4 I__11826 (
            .O(N__50011),
            .I(N__49998));
    LocalMux I__11825 (
            .O(N__50006),
            .I(N__49998));
    LocalMux I__11824 (
            .O(N__50003),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv12 I__11823 (
            .O(N__49998),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    CascadeMux I__11822 (
            .O(N__49993),
            .I(N__49990));
    InMux I__11821 (
            .O(N__49990),
            .I(N__49986));
    InMux I__11820 (
            .O(N__49989),
            .I(N__49983));
    LocalMux I__11819 (
            .O(N__49986),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    LocalMux I__11818 (
            .O(N__49983),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    ClkMux I__11817 (
            .O(N__49978),
            .I(N__49591));
    ClkMux I__11816 (
            .O(N__49977),
            .I(N__49591));
    ClkMux I__11815 (
            .O(N__49976),
            .I(N__49591));
    ClkMux I__11814 (
            .O(N__49975),
            .I(N__49591));
    ClkMux I__11813 (
            .O(N__49974),
            .I(N__49591));
    ClkMux I__11812 (
            .O(N__49973),
            .I(N__49591));
    ClkMux I__11811 (
            .O(N__49972),
            .I(N__49591));
    ClkMux I__11810 (
            .O(N__49971),
            .I(N__49591));
    ClkMux I__11809 (
            .O(N__49970),
            .I(N__49591));
    ClkMux I__11808 (
            .O(N__49969),
            .I(N__49591));
    ClkMux I__11807 (
            .O(N__49968),
            .I(N__49591));
    ClkMux I__11806 (
            .O(N__49967),
            .I(N__49591));
    ClkMux I__11805 (
            .O(N__49966),
            .I(N__49591));
    ClkMux I__11804 (
            .O(N__49965),
            .I(N__49591));
    ClkMux I__11803 (
            .O(N__49964),
            .I(N__49591));
    ClkMux I__11802 (
            .O(N__49963),
            .I(N__49591));
    ClkMux I__11801 (
            .O(N__49962),
            .I(N__49591));
    ClkMux I__11800 (
            .O(N__49961),
            .I(N__49591));
    ClkMux I__11799 (
            .O(N__49960),
            .I(N__49591));
    ClkMux I__11798 (
            .O(N__49959),
            .I(N__49591));
    ClkMux I__11797 (
            .O(N__49958),
            .I(N__49591));
    ClkMux I__11796 (
            .O(N__49957),
            .I(N__49591));
    ClkMux I__11795 (
            .O(N__49956),
            .I(N__49591));
    ClkMux I__11794 (
            .O(N__49955),
            .I(N__49591));
    ClkMux I__11793 (
            .O(N__49954),
            .I(N__49591));
    ClkMux I__11792 (
            .O(N__49953),
            .I(N__49591));
    ClkMux I__11791 (
            .O(N__49952),
            .I(N__49591));
    ClkMux I__11790 (
            .O(N__49951),
            .I(N__49591));
    ClkMux I__11789 (
            .O(N__49950),
            .I(N__49591));
    ClkMux I__11788 (
            .O(N__49949),
            .I(N__49591));
    ClkMux I__11787 (
            .O(N__49948),
            .I(N__49591));
    ClkMux I__11786 (
            .O(N__49947),
            .I(N__49591));
    ClkMux I__11785 (
            .O(N__49946),
            .I(N__49591));
    ClkMux I__11784 (
            .O(N__49945),
            .I(N__49591));
    ClkMux I__11783 (
            .O(N__49944),
            .I(N__49591));
    ClkMux I__11782 (
            .O(N__49943),
            .I(N__49591));
    ClkMux I__11781 (
            .O(N__49942),
            .I(N__49591));
    ClkMux I__11780 (
            .O(N__49941),
            .I(N__49591));
    ClkMux I__11779 (
            .O(N__49940),
            .I(N__49591));
    ClkMux I__11778 (
            .O(N__49939),
            .I(N__49591));
    ClkMux I__11777 (
            .O(N__49938),
            .I(N__49591));
    ClkMux I__11776 (
            .O(N__49937),
            .I(N__49591));
    ClkMux I__11775 (
            .O(N__49936),
            .I(N__49591));
    ClkMux I__11774 (
            .O(N__49935),
            .I(N__49591));
    ClkMux I__11773 (
            .O(N__49934),
            .I(N__49591));
    ClkMux I__11772 (
            .O(N__49933),
            .I(N__49591));
    ClkMux I__11771 (
            .O(N__49932),
            .I(N__49591));
    ClkMux I__11770 (
            .O(N__49931),
            .I(N__49591));
    ClkMux I__11769 (
            .O(N__49930),
            .I(N__49591));
    ClkMux I__11768 (
            .O(N__49929),
            .I(N__49591));
    ClkMux I__11767 (
            .O(N__49928),
            .I(N__49591));
    ClkMux I__11766 (
            .O(N__49927),
            .I(N__49591));
    ClkMux I__11765 (
            .O(N__49926),
            .I(N__49591));
    ClkMux I__11764 (
            .O(N__49925),
            .I(N__49591));
    ClkMux I__11763 (
            .O(N__49924),
            .I(N__49591));
    ClkMux I__11762 (
            .O(N__49923),
            .I(N__49591));
    ClkMux I__11761 (
            .O(N__49922),
            .I(N__49591));
    ClkMux I__11760 (
            .O(N__49921),
            .I(N__49591));
    ClkMux I__11759 (
            .O(N__49920),
            .I(N__49591));
    ClkMux I__11758 (
            .O(N__49919),
            .I(N__49591));
    ClkMux I__11757 (
            .O(N__49918),
            .I(N__49591));
    ClkMux I__11756 (
            .O(N__49917),
            .I(N__49591));
    ClkMux I__11755 (
            .O(N__49916),
            .I(N__49591));
    ClkMux I__11754 (
            .O(N__49915),
            .I(N__49591));
    ClkMux I__11753 (
            .O(N__49914),
            .I(N__49591));
    ClkMux I__11752 (
            .O(N__49913),
            .I(N__49591));
    ClkMux I__11751 (
            .O(N__49912),
            .I(N__49591));
    ClkMux I__11750 (
            .O(N__49911),
            .I(N__49591));
    ClkMux I__11749 (
            .O(N__49910),
            .I(N__49591));
    ClkMux I__11748 (
            .O(N__49909),
            .I(N__49591));
    ClkMux I__11747 (
            .O(N__49908),
            .I(N__49591));
    ClkMux I__11746 (
            .O(N__49907),
            .I(N__49591));
    ClkMux I__11745 (
            .O(N__49906),
            .I(N__49591));
    ClkMux I__11744 (
            .O(N__49905),
            .I(N__49591));
    ClkMux I__11743 (
            .O(N__49904),
            .I(N__49591));
    ClkMux I__11742 (
            .O(N__49903),
            .I(N__49591));
    ClkMux I__11741 (
            .O(N__49902),
            .I(N__49591));
    ClkMux I__11740 (
            .O(N__49901),
            .I(N__49591));
    ClkMux I__11739 (
            .O(N__49900),
            .I(N__49591));
    ClkMux I__11738 (
            .O(N__49899),
            .I(N__49591));
    ClkMux I__11737 (
            .O(N__49898),
            .I(N__49591));
    ClkMux I__11736 (
            .O(N__49897),
            .I(N__49591));
    ClkMux I__11735 (
            .O(N__49896),
            .I(N__49591));
    ClkMux I__11734 (
            .O(N__49895),
            .I(N__49591));
    ClkMux I__11733 (
            .O(N__49894),
            .I(N__49591));
    ClkMux I__11732 (
            .O(N__49893),
            .I(N__49591));
    ClkMux I__11731 (
            .O(N__49892),
            .I(N__49591));
    ClkMux I__11730 (
            .O(N__49891),
            .I(N__49591));
    ClkMux I__11729 (
            .O(N__49890),
            .I(N__49591));
    ClkMux I__11728 (
            .O(N__49889),
            .I(N__49591));
    ClkMux I__11727 (
            .O(N__49888),
            .I(N__49591));
    ClkMux I__11726 (
            .O(N__49887),
            .I(N__49591));
    ClkMux I__11725 (
            .O(N__49886),
            .I(N__49591));
    ClkMux I__11724 (
            .O(N__49885),
            .I(N__49591));
    ClkMux I__11723 (
            .O(N__49884),
            .I(N__49591));
    ClkMux I__11722 (
            .O(N__49883),
            .I(N__49591));
    ClkMux I__11721 (
            .O(N__49882),
            .I(N__49591));
    ClkMux I__11720 (
            .O(N__49881),
            .I(N__49591));
    ClkMux I__11719 (
            .O(N__49880),
            .I(N__49591));
    ClkMux I__11718 (
            .O(N__49879),
            .I(N__49591));
    ClkMux I__11717 (
            .O(N__49878),
            .I(N__49591));
    ClkMux I__11716 (
            .O(N__49877),
            .I(N__49591));
    ClkMux I__11715 (
            .O(N__49876),
            .I(N__49591));
    ClkMux I__11714 (
            .O(N__49875),
            .I(N__49591));
    ClkMux I__11713 (
            .O(N__49874),
            .I(N__49591));
    ClkMux I__11712 (
            .O(N__49873),
            .I(N__49591));
    ClkMux I__11711 (
            .O(N__49872),
            .I(N__49591));
    ClkMux I__11710 (
            .O(N__49871),
            .I(N__49591));
    ClkMux I__11709 (
            .O(N__49870),
            .I(N__49591));
    ClkMux I__11708 (
            .O(N__49869),
            .I(N__49591));
    ClkMux I__11707 (
            .O(N__49868),
            .I(N__49591));
    ClkMux I__11706 (
            .O(N__49867),
            .I(N__49591));
    ClkMux I__11705 (
            .O(N__49866),
            .I(N__49591));
    ClkMux I__11704 (
            .O(N__49865),
            .I(N__49591));
    ClkMux I__11703 (
            .O(N__49864),
            .I(N__49591));
    ClkMux I__11702 (
            .O(N__49863),
            .I(N__49591));
    ClkMux I__11701 (
            .O(N__49862),
            .I(N__49591));
    ClkMux I__11700 (
            .O(N__49861),
            .I(N__49591));
    ClkMux I__11699 (
            .O(N__49860),
            .I(N__49591));
    ClkMux I__11698 (
            .O(N__49859),
            .I(N__49591));
    ClkMux I__11697 (
            .O(N__49858),
            .I(N__49591));
    ClkMux I__11696 (
            .O(N__49857),
            .I(N__49591));
    ClkMux I__11695 (
            .O(N__49856),
            .I(N__49591));
    ClkMux I__11694 (
            .O(N__49855),
            .I(N__49591));
    ClkMux I__11693 (
            .O(N__49854),
            .I(N__49591));
    ClkMux I__11692 (
            .O(N__49853),
            .I(N__49591));
    ClkMux I__11691 (
            .O(N__49852),
            .I(N__49591));
    ClkMux I__11690 (
            .O(N__49851),
            .I(N__49591));
    ClkMux I__11689 (
            .O(N__49850),
            .I(N__49591));
    GlobalMux I__11688 (
            .O(N__49591),
            .I(clk_100mhz_0));
    InMux I__11687 (
            .O(N__49588),
            .I(N__49577));
    InMux I__11686 (
            .O(N__49587),
            .I(N__49574));
    InMux I__11685 (
            .O(N__49586),
            .I(N__49571));
    InMux I__11684 (
            .O(N__49585),
            .I(N__49568));
    InMux I__11683 (
            .O(N__49584),
            .I(N__49565));
    InMux I__11682 (
            .O(N__49583),
            .I(N__49562));
    InMux I__11681 (
            .O(N__49582),
            .I(N__49559));
    InMux I__11680 (
            .O(N__49581),
            .I(N__49554));
    InMux I__11679 (
            .O(N__49580),
            .I(N__49554));
    LocalMux I__11678 (
            .O(N__49577),
            .I(N__49551));
    LocalMux I__11677 (
            .O(N__49574),
            .I(N__49548));
    LocalMux I__11676 (
            .O(N__49571),
            .I(N__49545));
    LocalMux I__11675 (
            .O(N__49568),
            .I(N__49475));
    LocalMux I__11674 (
            .O(N__49565),
            .I(N__49453));
    LocalMux I__11673 (
            .O(N__49562),
            .I(N__49445));
    LocalMux I__11672 (
            .O(N__49559),
            .I(N__49427));
    LocalMux I__11671 (
            .O(N__49554),
            .I(N__49417));
    Glb2LocalMux I__11670 (
            .O(N__49551),
            .I(N__49138));
    Glb2LocalMux I__11669 (
            .O(N__49548),
            .I(N__49138));
    Glb2LocalMux I__11668 (
            .O(N__49545),
            .I(N__49138));
    SRMux I__11667 (
            .O(N__49544),
            .I(N__49138));
    SRMux I__11666 (
            .O(N__49543),
            .I(N__49138));
    SRMux I__11665 (
            .O(N__49542),
            .I(N__49138));
    SRMux I__11664 (
            .O(N__49541),
            .I(N__49138));
    SRMux I__11663 (
            .O(N__49540),
            .I(N__49138));
    SRMux I__11662 (
            .O(N__49539),
            .I(N__49138));
    SRMux I__11661 (
            .O(N__49538),
            .I(N__49138));
    SRMux I__11660 (
            .O(N__49537),
            .I(N__49138));
    SRMux I__11659 (
            .O(N__49536),
            .I(N__49138));
    SRMux I__11658 (
            .O(N__49535),
            .I(N__49138));
    SRMux I__11657 (
            .O(N__49534),
            .I(N__49138));
    SRMux I__11656 (
            .O(N__49533),
            .I(N__49138));
    SRMux I__11655 (
            .O(N__49532),
            .I(N__49138));
    SRMux I__11654 (
            .O(N__49531),
            .I(N__49138));
    SRMux I__11653 (
            .O(N__49530),
            .I(N__49138));
    SRMux I__11652 (
            .O(N__49529),
            .I(N__49138));
    SRMux I__11651 (
            .O(N__49528),
            .I(N__49138));
    SRMux I__11650 (
            .O(N__49527),
            .I(N__49138));
    SRMux I__11649 (
            .O(N__49526),
            .I(N__49138));
    SRMux I__11648 (
            .O(N__49525),
            .I(N__49138));
    SRMux I__11647 (
            .O(N__49524),
            .I(N__49138));
    SRMux I__11646 (
            .O(N__49523),
            .I(N__49138));
    SRMux I__11645 (
            .O(N__49522),
            .I(N__49138));
    SRMux I__11644 (
            .O(N__49521),
            .I(N__49138));
    SRMux I__11643 (
            .O(N__49520),
            .I(N__49138));
    SRMux I__11642 (
            .O(N__49519),
            .I(N__49138));
    SRMux I__11641 (
            .O(N__49518),
            .I(N__49138));
    SRMux I__11640 (
            .O(N__49517),
            .I(N__49138));
    SRMux I__11639 (
            .O(N__49516),
            .I(N__49138));
    SRMux I__11638 (
            .O(N__49515),
            .I(N__49138));
    SRMux I__11637 (
            .O(N__49514),
            .I(N__49138));
    SRMux I__11636 (
            .O(N__49513),
            .I(N__49138));
    SRMux I__11635 (
            .O(N__49512),
            .I(N__49138));
    SRMux I__11634 (
            .O(N__49511),
            .I(N__49138));
    SRMux I__11633 (
            .O(N__49510),
            .I(N__49138));
    SRMux I__11632 (
            .O(N__49509),
            .I(N__49138));
    SRMux I__11631 (
            .O(N__49508),
            .I(N__49138));
    SRMux I__11630 (
            .O(N__49507),
            .I(N__49138));
    SRMux I__11629 (
            .O(N__49506),
            .I(N__49138));
    SRMux I__11628 (
            .O(N__49505),
            .I(N__49138));
    SRMux I__11627 (
            .O(N__49504),
            .I(N__49138));
    SRMux I__11626 (
            .O(N__49503),
            .I(N__49138));
    SRMux I__11625 (
            .O(N__49502),
            .I(N__49138));
    SRMux I__11624 (
            .O(N__49501),
            .I(N__49138));
    SRMux I__11623 (
            .O(N__49500),
            .I(N__49138));
    SRMux I__11622 (
            .O(N__49499),
            .I(N__49138));
    SRMux I__11621 (
            .O(N__49498),
            .I(N__49138));
    SRMux I__11620 (
            .O(N__49497),
            .I(N__49138));
    SRMux I__11619 (
            .O(N__49496),
            .I(N__49138));
    SRMux I__11618 (
            .O(N__49495),
            .I(N__49138));
    SRMux I__11617 (
            .O(N__49494),
            .I(N__49138));
    SRMux I__11616 (
            .O(N__49493),
            .I(N__49138));
    SRMux I__11615 (
            .O(N__49492),
            .I(N__49138));
    SRMux I__11614 (
            .O(N__49491),
            .I(N__49138));
    SRMux I__11613 (
            .O(N__49490),
            .I(N__49138));
    SRMux I__11612 (
            .O(N__49489),
            .I(N__49138));
    SRMux I__11611 (
            .O(N__49488),
            .I(N__49138));
    SRMux I__11610 (
            .O(N__49487),
            .I(N__49138));
    SRMux I__11609 (
            .O(N__49486),
            .I(N__49138));
    SRMux I__11608 (
            .O(N__49485),
            .I(N__49138));
    SRMux I__11607 (
            .O(N__49484),
            .I(N__49138));
    SRMux I__11606 (
            .O(N__49483),
            .I(N__49138));
    SRMux I__11605 (
            .O(N__49482),
            .I(N__49138));
    SRMux I__11604 (
            .O(N__49481),
            .I(N__49138));
    SRMux I__11603 (
            .O(N__49480),
            .I(N__49138));
    SRMux I__11602 (
            .O(N__49479),
            .I(N__49138));
    SRMux I__11601 (
            .O(N__49478),
            .I(N__49138));
    Glb2LocalMux I__11600 (
            .O(N__49475),
            .I(N__49138));
    SRMux I__11599 (
            .O(N__49474),
            .I(N__49138));
    SRMux I__11598 (
            .O(N__49473),
            .I(N__49138));
    SRMux I__11597 (
            .O(N__49472),
            .I(N__49138));
    SRMux I__11596 (
            .O(N__49471),
            .I(N__49138));
    SRMux I__11595 (
            .O(N__49470),
            .I(N__49138));
    SRMux I__11594 (
            .O(N__49469),
            .I(N__49138));
    SRMux I__11593 (
            .O(N__49468),
            .I(N__49138));
    SRMux I__11592 (
            .O(N__49467),
            .I(N__49138));
    SRMux I__11591 (
            .O(N__49466),
            .I(N__49138));
    SRMux I__11590 (
            .O(N__49465),
            .I(N__49138));
    SRMux I__11589 (
            .O(N__49464),
            .I(N__49138));
    SRMux I__11588 (
            .O(N__49463),
            .I(N__49138));
    SRMux I__11587 (
            .O(N__49462),
            .I(N__49138));
    SRMux I__11586 (
            .O(N__49461),
            .I(N__49138));
    SRMux I__11585 (
            .O(N__49460),
            .I(N__49138));
    SRMux I__11584 (
            .O(N__49459),
            .I(N__49138));
    SRMux I__11583 (
            .O(N__49458),
            .I(N__49138));
    SRMux I__11582 (
            .O(N__49457),
            .I(N__49138));
    SRMux I__11581 (
            .O(N__49456),
            .I(N__49138));
    Glb2LocalMux I__11580 (
            .O(N__49453),
            .I(N__49138));
    SRMux I__11579 (
            .O(N__49452),
            .I(N__49138));
    SRMux I__11578 (
            .O(N__49451),
            .I(N__49138));
    SRMux I__11577 (
            .O(N__49450),
            .I(N__49138));
    SRMux I__11576 (
            .O(N__49449),
            .I(N__49138));
    SRMux I__11575 (
            .O(N__49448),
            .I(N__49138));
    Glb2LocalMux I__11574 (
            .O(N__49445),
            .I(N__49138));
    SRMux I__11573 (
            .O(N__49444),
            .I(N__49138));
    SRMux I__11572 (
            .O(N__49443),
            .I(N__49138));
    SRMux I__11571 (
            .O(N__49442),
            .I(N__49138));
    SRMux I__11570 (
            .O(N__49441),
            .I(N__49138));
    SRMux I__11569 (
            .O(N__49440),
            .I(N__49138));
    SRMux I__11568 (
            .O(N__49439),
            .I(N__49138));
    SRMux I__11567 (
            .O(N__49438),
            .I(N__49138));
    SRMux I__11566 (
            .O(N__49437),
            .I(N__49138));
    SRMux I__11565 (
            .O(N__49436),
            .I(N__49138));
    SRMux I__11564 (
            .O(N__49435),
            .I(N__49138));
    SRMux I__11563 (
            .O(N__49434),
            .I(N__49138));
    SRMux I__11562 (
            .O(N__49433),
            .I(N__49138));
    SRMux I__11561 (
            .O(N__49432),
            .I(N__49138));
    SRMux I__11560 (
            .O(N__49431),
            .I(N__49138));
    SRMux I__11559 (
            .O(N__49430),
            .I(N__49138));
    Glb2LocalMux I__11558 (
            .O(N__49427),
            .I(N__49138));
    SRMux I__11557 (
            .O(N__49426),
            .I(N__49138));
    SRMux I__11556 (
            .O(N__49425),
            .I(N__49138));
    SRMux I__11555 (
            .O(N__49424),
            .I(N__49138));
    SRMux I__11554 (
            .O(N__49423),
            .I(N__49138));
    SRMux I__11553 (
            .O(N__49422),
            .I(N__49138));
    SRMux I__11552 (
            .O(N__49421),
            .I(N__49138));
    SRMux I__11551 (
            .O(N__49420),
            .I(N__49138));
    Glb2LocalMux I__11550 (
            .O(N__49417),
            .I(N__49138));
    SRMux I__11549 (
            .O(N__49416),
            .I(N__49138));
    SRMux I__11548 (
            .O(N__49415),
            .I(N__49138));
    SRMux I__11547 (
            .O(N__49414),
            .I(N__49138));
    SRMux I__11546 (
            .O(N__49413),
            .I(N__49138));
    SRMux I__11545 (
            .O(N__49412),
            .I(N__49138));
    SRMux I__11544 (
            .O(N__49411),
            .I(N__49138));
    SRMux I__11543 (
            .O(N__49410),
            .I(N__49138));
    SRMux I__11542 (
            .O(N__49409),
            .I(N__49138));
    SRMux I__11541 (
            .O(N__49408),
            .I(N__49138));
    SRMux I__11540 (
            .O(N__49407),
            .I(N__49138));
    SRMux I__11539 (
            .O(N__49406),
            .I(N__49138));
    SRMux I__11538 (
            .O(N__49405),
            .I(N__49138));
    GlobalMux I__11537 (
            .O(N__49138),
            .I(N__49135));
    gio2CtrlBuf I__11536 (
            .O(N__49135),
            .I(red_c_g));
    InMux I__11535 (
            .O(N__49132),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__11534 (
            .O(N__49129),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__11533 (
            .O(N__49126),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    CEMux I__11532 (
            .O(N__49123),
            .I(N__49117));
    CEMux I__11531 (
            .O(N__49122),
            .I(N__49114));
    CEMux I__11530 (
            .O(N__49121),
            .I(N__49111));
    CEMux I__11529 (
            .O(N__49120),
            .I(N__49105));
    LocalMux I__11528 (
            .O(N__49117),
            .I(N__49095));
    LocalMux I__11527 (
            .O(N__49114),
            .I(N__49076));
    LocalMux I__11526 (
            .O(N__49111),
            .I(N__49073));
    CEMux I__11525 (
            .O(N__49110),
            .I(N__49070));
    CEMux I__11524 (
            .O(N__49109),
            .I(N__49066));
    CEMux I__11523 (
            .O(N__49108),
            .I(N__49063));
    LocalMux I__11522 (
            .O(N__49105),
            .I(N__49060));
    InMux I__11521 (
            .O(N__49104),
            .I(N__49051));
    InMux I__11520 (
            .O(N__49103),
            .I(N__49051));
    InMux I__11519 (
            .O(N__49102),
            .I(N__49051));
    InMux I__11518 (
            .O(N__49101),
            .I(N__49051));
    InMux I__11517 (
            .O(N__49100),
            .I(N__49044));
    InMux I__11516 (
            .O(N__49099),
            .I(N__49044));
    InMux I__11515 (
            .O(N__49098),
            .I(N__49044));
    Span4Mux_h I__11514 (
            .O(N__49095),
            .I(N__49041));
    InMux I__11513 (
            .O(N__49094),
            .I(N__49032));
    InMux I__11512 (
            .O(N__49093),
            .I(N__49032));
    InMux I__11511 (
            .O(N__49092),
            .I(N__49032));
    InMux I__11510 (
            .O(N__49091),
            .I(N__49032));
    InMux I__11509 (
            .O(N__49090),
            .I(N__49023));
    InMux I__11508 (
            .O(N__49089),
            .I(N__49023));
    InMux I__11507 (
            .O(N__49088),
            .I(N__49023));
    InMux I__11506 (
            .O(N__49087),
            .I(N__49023));
    InMux I__11505 (
            .O(N__49086),
            .I(N__49014));
    InMux I__11504 (
            .O(N__49085),
            .I(N__49014));
    InMux I__11503 (
            .O(N__49084),
            .I(N__49014));
    InMux I__11502 (
            .O(N__49083),
            .I(N__49014));
    InMux I__11501 (
            .O(N__49082),
            .I(N__49005));
    InMux I__11500 (
            .O(N__49081),
            .I(N__49005));
    InMux I__11499 (
            .O(N__49080),
            .I(N__49005));
    InMux I__11498 (
            .O(N__49079),
            .I(N__49005));
    Span4Mux_h I__11497 (
            .O(N__49076),
            .I(N__48998));
    Span4Mux_h I__11496 (
            .O(N__49073),
            .I(N__48998));
    LocalMux I__11495 (
            .O(N__49070),
            .I(N__48998));
    CEMux I__11494 (
            .O(N__49069),
            .I(N__48995));
    LocalMux I__11493 (
            .O(N__49066),
            .I(N__48990));
    LocalMux I__11492 (
            .O(N__49063),
            .I(N__48987));
    Span4Mux_v I__11491 (
            .O(N__49060),
            .I(N__48980));
    LocalMux I__11490 (
            .O(N__49051),
            .I(N__48975));
    LocalMux I__11489 (
            .O(N__49044),
            .I(N__48975));
    Span4Mux_h I__11488 (
            .O(N__49041),
            .I(N__48964));
    LocalMux I__11487 (
            .O(N__49032),
            .I(N__48964));
    LocalMux I__11486 (
            .O(N__49023),
            .I(N__48964));
    LocalMux I__11485 (
            .O(N__49014),
            .I(N__48964));
    LocalMux I__11484 (
            .O(N__49005),
            .I(N__48964));
    Span4Mux_v I__11483 (
            .O(N__48998),
            .I(N__48958));
    LocalMux I__11482 (
            .O(N__48995),
            .I(N__48955));
    InMux I__11481 (
            .O(N__48994),
            .I(N__48952));
    CEMux I__11480 (
            .O(N__48993),
            .I(N__48948));
    Span12Mux_h I__11479 (
            .O(N__48990),
            .I(N__48943));
    Sp12to4 I__11478 (
            .O(N__48987),
            .I(N__48943));
    InMux I__11477 (
            .O(N__48986),
            .I(N__48934));
    InMux I__11476 (
            .O(N__48985),
            .I(N__48934));
    InMux I__11475 (
            .O(N__48984),
            .I(N__48934));
    InMux I__11474 (
            .O(N__48983),
            .I(N__48934));
    Span4Mux_h I__11473 (
            .O(N__48980),
            .I(N__48929));
    Span4Mux_v I__11472 (
            .O(N__48975),
            .I(N__48929));
    Span4Mux_v I__11471 (
            .O(N__48964),
            .I(N__48926));
    InMux I__11470 (
            .O(N__48963),
            .I(N__48919));
    InMux I__11469 (
            .O(N__48962),
            .I(N__48919));
    InMux I__11468 (
            .O(N__48961),
            .I(N__48919));
    Span4Mux_h I__11467 (
            .O(N__48958),
            .I(N__48912));
    Span4Mux_v I__11466 (
            .O(N__48955),
            .I(N__48912));
    LocalMux I__11465 (
            .O(N__48952),
            .I(N__48912));
    CEMux I__11464 (
            .O(N__48951),
            .I(N__48909));
    LocalMux I__11463 (
            .O(N__48948),
            .I(N__48896));
    Span12Mux_v I__11462 (
            .O(N__48943),
            .I(N__48896));
    LocalMux I__11461 (
            .O(N__48934),
            .I(N__48896));
    Sp12to4 I__11460 (
            .O(N__48929),
            .I(N__48896));
    Sp12to4 I__11459 (
            .O(N__48926),
            .I(N__48896));
    LocalMux I__11458 (
            .O(N__48919),
            .I(N__48896));
    Span4Mux_v I__11457 (
            .O(N__48912),
            .I(N__48893));
    LocalMux I__11456 (
            .O(N__48909),
            .I(N__48888));
    Span12Mux_s9_h I__11455 (
            .O(N__48896),
            .I(N__48888));
    Odrv4 I__11454 (
            .O(N__48893),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__11453 (
            .O(N__48888),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__11452 (
            .O(N__48883),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__11451 (
            .O(N__48880),
            .I(N__48877));
    LocalMux I__11450 (
            .O(N__48877),
            .I(N__48873));
    InMux I__11449 (
            .O(N__48876),
            .I(N__48870));
    Span4Mux_v I__11448 (
            .O(N__48873),
            .I(N__48867));
    LocalMux I__11447 (
            .O(N__48870),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__11446 (
            .O(N__48867),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__11445 (
            .O(N__48862),
            .I(N__48858));
    InMux I__11444 (
            .O(N__48861),
            .I(N__48855));
    LocalMux I__11443 (
            .O(N__48858),
            .I(N__48852));
    LocalMux I__11442 (
            .O(N__48855),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv12 I__11441 (
            .O(N__48852),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__11440 (
            .O(N__48847),
            .I(N__48844));
    LocalMux I__11439 (
            .O(N__48844),
            .I(N__48841));
    Span4Mux_h I__11438 (
            .O(N__48841),
            .I(N__48838));
    Span4Mux_v I__11437 (
            .O(N__48838),
            .I(N__48835));
    Odrv4 I__11436 (
            .O(N__48835),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df20 ));
    InMux I__11435 (
            .O(N__48832),
            .I(N__48828));
    InMux I__11434 (
            .O(N__48831),
            .I(N__48825));
    LocalMux I__11433 (
            .O(N__48828),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__11432 (
            .O(N__48825),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__11431 (
            .O(N__48820),
            .I(N__48816));
    InMux I__11430 (
            .O(N__48819),
            .I(N__48813));
    LocalMux I__11429 (
            .O(N__48816),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__11428 (
            .O(N__48813),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__11427 (
            .O(N__48808),
            .I(N__48805));
    LocalMux I__11426 (
            .O(N__48805),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df26 ));
    InMux I__11425 (
            .O(N__48802),
            .I(N__48798));
    InMux I__11424 (
            .O(N__48801),
            .I(N__48795));
    LocalMux I__11423 (
            .O(N__48798),
            .I(N__48792));
    LocalMux I__11422 (
            .O(N__48795),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__11421 (
            .O(N__48792),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__11420 (
            .O(N__48787),
            .I(N__48783));
    InMux I__11419 (
            .O(N__48786),
            .I(N__48780));
    LocalMux I__11418 (
            .O(N__48783),
            .I(N__48777));
    LocalMux I__11417 (
            .O(N__48780),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__11416 (
            .O(N__48777),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__11415 (
            .O(N__48772),
            .I(N__48769));
    LocalMux I__11414 (
            .O(N__48769),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df22 ));
    InMux I__11413 (
            .O(N__48766),
            .I(N__48762));
    InMux I__11412 (
            .O(N__48765),
            .I(N__48759));
    LocalMux I__11411 (
            .O(N__48762),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__11410 (
            .O(N__48759),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__11409 (
            .O(N__48754),
            .I(N__48750));
    InMux I__11408 (
            .O(N__48753),
            .I(N__48747));
    LocalMux I__11407 (
            .O(N__48750),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__11406 (
            .O(N__48747),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__11405 (
            .O(N__48742),
            .I(N__48739));
    LocalMux I__11404 (
            .O(N__48739),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df28 ));
    InMux I__11403 (
            .O(N__48736),
            .I(N__48731));
    InMux I__11402 (
            .O(N__48735),
            .I(N__48728));
    InMux I__11401 (
            .O(N__48734),
            .I(N__48725));
    LocalMux I__11400 (
            .O(N__48731),
            .I(N__48722));
    LocalMux I__11399 (
            .O(N__48728),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__11398 (
            .O(N__48725),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__11397 (
            .O(N__48722),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    CascadeMux I__11396 (
            .O(N__48715),
            .I(N__48712));
    InMux I__11395 (
            .O(N__48712),
            .I(N__48707));
    CascadeMux I__11394 (
            .O(N__48711),
            .I(N__48703));
    InMux I__11393 (
            .O(N__48710),
            .I(N__48700));
    LocalMux I__11392 (
            .O(N__48707),
            .I(N__48697));
    InMux I__11391 (
            .O(N__48706),
            .I(N__48694));
    InMux I__11390 (
            .O(N__48703),
            .I(N__48691));
    LocalMux I__11389 (
            .O(N__48700),
            .I(N__48686));
    Span4Mux_h I__11388 (
            .O(N__48697),
            .I(N__48686));
    LocalMux I__11387 (
            .O(N__48694),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    LocalMux I__11386 (
            .O(N__48691),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__11385 (
            .O(N__48686),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__11384 (
            .O(N__48679),
            .I(N__48676));
    LocalMux I__11383 (
            .O(N__48676),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    CascadeMux I__11382 (
            .O(N__48673),
            .I(N__48670));
    InMux I__11381 (
            .O(N__48670),
            .I(N__48666));
    InMux I__11380 (
            .O(N__48669),
            .I(N__48662));
    LocalMux I__11379 (
            .O(N__48666),
            .I(N__48659));
    InMux I__11378 (
            .O(N__48665),
            .I(N__48656));
    LocalMux I__11377 (
            .O(N__48662),
            .I(N__48651));
    Span4Mux_v I__11376 (
            .O(N__48659),
            .I(N__48651));
    LocalMux I__11375 (
            .O(N__48656),
            .I(N__48648));
    Odrv4 I__11374 (
            .O(N__48651),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__11373 (
            .O(N__48648),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__11372 (
            .O(N__48643),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__11371 (
            .O(N__48640),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__11370 (
            .O(N__48637),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__11369 (
            .O(N__48634),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__11368 (
            .O(N__48631),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__11367 (
            .O(N__48628),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__11366 (
            .O(N__48625),
            .I(bfn_18_20_0_));
    InMux I__11365 (
            .O(N__48622),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__11364 (
            .O(N__48619),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__11363 (
            .O(N__48616),
            .I(N__48612));
    InMux I__11362 (
            .O(N__48615),
            .I(N__48609));
    LocalMux I__11361 (
            .O(N__48612),
            .I(N__48606));
    LocalMux I__11360 (
            .O(N__48609),
            .I(N__48601));
    Span4Mux_v I__11359 (
            .O(N__48606),
            .I(N__48601));
    Odrv4 I__11358 (
            .O(N__48601),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__11357 (
            .O(N__48598),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__11356 (
            .O(N__48595),
            .I(N__48591));
    InMux I__11355 (
            .O(N__48594),
            .I(N__48588));
    LocalMux I__11354 (
            .O(N__48591),
            .I(N__48585));
    LocalMux I__11353 (
            .O(N__48588),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__11352 (
            .O(N__48585),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__11351 (
            .O(N__48580),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__11350 (
            .O(N__48577),
            .I(N__48573));
    InMux I__11349 (
            .O(N__48576),
            .I(N__48570));
    LocalMux I__11348 (
            .O(N__48573),
            .I(N__48567));
    LocalMux I__11347 (
            .O(N__48570),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__11346 (
            .O(N__48567),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__11345 (
            .O(N__48562),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__11344 (
            .O(N__48559),
            .I(N__48555));
    InMux I__11343 (
            .O(N__48558),
            .I(N__48552));
    LocalMux I__11342 (
            .O(N__48555),
            .I(N__48549));
    LocalMux I__11341 (
            .O(N__48552),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__11340 (
            .O(N__48549),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__11339 (
            .O(N__48544),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__11338 (
            .O(N__48541),
            .I(N__48537));
    InMux I__11337 (
            .O(N__48540),
            .I(N__48534));
    LocalMux I__11336 (
            .O(N__48537),
            .I(N__48531));
    LocalMux I__11335 (
            .O(N__48534),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__11334 (
            .O(N__48531),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__11333 (
            .O(N__48526),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    CascadeMux I__11332 (
            .O(N__48523),
            .I(N__48520));
    InMux I__11331 (
            .O(N__48520),
            .I(N__48514));
    InMux I__11330 (
            .O(N__48519),
            .I(N__48514));
    LocalMux I__11329 (
            .O(N__48514),
            .I(N__48510));
    InMux I__11328 (
            .O(N__48513),
            .I(N__48507));
    Span4Mux_h I__11327 (
            .O(N__48510),
            .I(N__48504));
    LocalMux I__11326 (
            .O(N__48507),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__11325 (
            .O(N__48504),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__11324 (
            .O(N__48499),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__11323 (
            .O(N__48496),
            .I(N__48489));
    InMux I__11322 (
            .O(N__48495),
            .I(N__48489));
    InMux I__11321 (
            .O(N__48494),
            .I(N__48486));
    LocalMux I__11320 (
            .O(N__48489),
            .I(N__48483));
    LocalMux I__11319 (
            .O(N__48486),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__11318 (
            .O(N__48483),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__11317 (
            .O(N__48478),
            .I(bfn_18_19_0_));
    CascadeMux I__11316 (
            .O(N__48475),
            .I(N__48471));
    InMux I__11315 (
            .O(N__48474),
            .I(N__48468));
    InMux I__11314 (
            .O(N__48471),
            .I(N__48464));
    LocalMux I__11313 (
            .O(N__48468),
            .I(N__48461));
    InMux I__11312 (
            .O(N__48467),
            .I(N__48458));
    LocalMux I__11311 (
            .O(N__48464),
            .I(N__48455));
    Span4Mux_h I__11310 (
            .O(N__48461),
            .I(N__48452));
    LocalMux I__11309 (
            .O(N__48458),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv12 I__11308 (
            .O(N__48455),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__11307 (
            .O(N__48452),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__11306 (
            .O(N__48445),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__11305 (
            .O(N__48442),
            .I(N__48439));
    LocalMux I__11304 (
            .O(N__48439),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28 ));
    CascadeMux I__11303 (
            .O(N__48436),
            .I(N__48432));
    InMux I__11302 (
            .O(N__48435),
            .I(N__48429));
    InMux I__11301 (
            .O(N__48432),
            .I(N__48426));
    LocalMux I__11300 (
            .O(N__48429),
            .I(N__48423));
    LocalMux I__11299 (
            .O(N__48426),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__11298 (
            .O(N__48423),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__11297 (
            .O(N__48418),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__11296 (
            .O(N__48415),
            .I(N__48411));
    InMux I__11295 (
            .O(N__48414),
            .I(N__48408));
    LocalMux I__11294 (
            .O(N__48411),
            .I(N__48405));
    LocalMux I__11293 (
            .O(N__48408),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__11292 (
            .O(N__48405),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__11291 (
            .O(N__48400),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__11290 (
            .O(N__48397),
            .I(N__48393));
    InMux I__11289 (
            .O(N__48396),
            .I(N__48390));
    LocalMux I__11288 (
            .O(N__48393),
            .I(N__48387));
    LocalMux I__11287 (
            .O(N__48390),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__11286 (
            .O(N__48387),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__11285 (
            .O(N__48382),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__11284 (
            .O(N__48379),
            .I(N__48375));
    InMux I__11283 (
            .O(N__48378),
            .I(N__48372));
    LocalMux I__11282 (
            .O(N__48375),
            .I(N__48369));
    LocalMux I__11281 (
            .O(N__48372),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__11280 (
            .O(N__48369),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__11279 (
            .O(N__48364),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__11278 (
            .O(N__48361),
            .I(N__48357));
    InMux I__11277 (
            .O(N__48360),
            .I(N__48354));
    LocalMux I__11276 (
            .O(N__48357),
            .I(N__48351));
    LocalMux I__11275 (
            .O(N__48354),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__11274 (
            .O(N__48351),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__11273 (
            .O(N__48346),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__11272 (
            .O(N__48343),
            .I(N__48339));
    InMux I__11271 (
            .O(N__48342),
            .I(N__48336));
    LocalMux I__11270 (
            .O(N__48339),
            .I(N__48333));
    LocalMux I__11269 (
            .O(N__48336),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__11268 (
            .O(N__48333),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__11267 (
            .O(N__48328),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__11266 (
            .O(N__48325),
            .I(N__48321));
    InMux I__11265 (
            .O(N__48324),
            .I(N__48318));
    LocalMux I__11264 (
            .O(N__48321),
            .I(N__48315));
    LocalMux I__11263 (
            .O(N__48318),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__11262 (
            .O(N__48315),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__11261 (
            .O(N__48310),
            .I(bfn_18_18_0_));
    InMux I__11260 (
            .O(N__48307),
            .I(N__48304));
    LocalMux I__11259 (
            .O(N__48304),
            .I(N__48300));
    InMux I__11258 (
            .O(N__48303),
            .I(N__48297));
    Span4Mux_v I__11257 (
            .O(N__48300),
            .I(N__48294));
    LocalMux I__11256 (
            .O(N__48297),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__11255 (
            .O(N__48294),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__11254 (
            .O(N__48289),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__11253 (
            .O(N__48286),
            .I(N__48283));
    LocalMux I__11252 (
            .O(N__48283),
            .I(N__48280));
    Span4Mux_v I__11251 (
            .O(N__48280),
            .I(N__48276));
    InMux I__11250 (
            .O(N__48279),
            .I(N__48273));
    Span4Mux_h I__11249 (
            .O(N__48276),
            .I(N__48270));
    LocalMux I__11248 (
            .O(N__48273),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__11247 (
            .O(N__48270),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__11246 (
            .O(N__48265),
            .I(bfn_18_16_0_));
    InMux I__11245 (
            .O(N__48262),
            .I(N__48258));
    InMux I__11244 (
            .O(N__48261),
            .I(N__48255));
    LocalMux I__11243 (
            .O(N__48258),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__11242 (
            .O(N__48255),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__11241 (
            .O(N__48250),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__11240 (
            .O(N__48247),
            .I(N__48243));
    InMux I__11239 (
            .O(N__48246),
            .I(N__48240));
    LocalMux I__11238 (
            .O(N__48243),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__11237 (
            .O(N__48240),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__11236 (
            .O(N__48235),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__11235 (
            .O(N__48232),
            .I(N__48228));
    InMux I__11234 (
            .O(N__48231),
            .I(N__48225));
    LocalMux I__11233 (
            .O(N__48228),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    LocalMux I__11232 (
            .O(N__48225),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__11231 (
            .O(N__48220),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__11230 (
            .O(N__48217),
            .I(N__48213));
    InMux I__11229 (
            .O(N__48216),
            .I(N__48210));
    LocalMux I__11228 (
            .O(N__48213),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    LocalMux I__11227 (
            .O(N__48210),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__11226 (
            .O(N__48205),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__11225 (
            .O(N__48202),
            .I(N__48197));
    InMux I__11224 (
            .O(N__48201),
            .I(N__48194));
    InMux I__11223 (
            .O(N__48200),
            .I(N__48191));
    LocalMux I__11222 (
            .O(N__48197),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__11221 (
            .O(N__48194),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    LocalMux I__11220 (
            .O(N__48191),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__11219 (
            .O(N__48184),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__11218 (
            .O(N__48181),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    CascadeMux I__11217 (
            .O(N__48178),
            .I(N__48175));
    InMux I__11216 (
            .O(N__48175),
            .I(N__48172));
    LocalMux I__11215 (
            .O(N__48172),
            .I(N__48167));
    CascadeMux I__11214 (
            .O(N__48171),
            .I(N__48163));
    InMux I__11213 (
            .O(N__48170),
            .I(N__48160));
    Span4Mux_h I__11212 (
            .O(N__48167),
            .I(N__48157));
    InMux I__11211 (
            .O(N__48166),
            .I(N__48154));
    InMux I__11210 (
            .O(N__48163),
            .I(N__48151));
    LocalMux I__11209 (
            .O(N__48160),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__11208 (
            .O(N__48157),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__11207 (
            .O(N__48154),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    LocalMux I__11206 (
            .O(N__48151),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__11205 (
            .O(N__48142),
            .I(N__48137));
    InMux I__11204 (
            .O(N__48141),
            .I(N__48134));
    InMux I__11203 (
            .O(N__48140),
            .I(N__48131));
    LocalMux I__11202 (
            .O(N__48137),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__11201 (
            .O(N__48134),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__11200 (
            .O(N__48131),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__11199 (
            .O(N__48124),
            .I(N__48121));
    InMux I__11198 (
            .O(N__48121),
            .I(N__48118));
    LocalMux I__11197 (
            .O(N__48118),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    InMux I__11196 (
            .O(N__48115),
            .I(N__48111));
    InMux I__11195 (
            .O(N__48114),
            .I(N__48108));
    LocalMux I__11194 (
            .O(N__48111),
            .I(N__48105));
    LocalMux I__11193 (
            .O(N__48108),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__11192 (
            .O(N__48105),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__11191 (
            .O(N__48100),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__11190 (
            .O(N__48097),
            .I(N__48094));
    InMux I__11189 (
            .O(N__48094),
            .I(N__48088));
    InMux I__11188 (
            .O(N__48093),
            .I(N__48088));
    LocalMux I__11187 (
            .O(N__48088),
            .I(N__48084));
    InMux I__11186 (
            .O(N__48087),
            .I(N__48081));
    Span4Mux_v I__11185 (
            .O(N__48084),
            .I(N__48078));
    LocalMux I__11184 (
            .O(N__48081),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__11183 (
            .O(N__48078),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__11182 (
            .O(N__48073),
            .I(bfn_18_15_0_));
    InMux I__11181 (
            .O(N__48070),
            .I(N__48064));
    InMux I__11180 (
            .O(N__48069),
            .I(N__48064));
    LocalMux I__11179 (
            .O(N__48064),
            .I(N__48060));
    InMux I__11178 (
            .O(N__48063),
            .I(N__48057));
    Span4Mux_v I__11177 (
            .O(N__48060),
            .I(N__48054));
    LocalMux I__11176 (
            .O(N__48057),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__11175 (
            .O(N__48054),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__11174 (
            .O(N__48049),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    CascadeMux I__11173 (
            .O(N__48046),
            .I(N__48043));
    InMux I__11172 (
            .O(N__48043),
            .I(N__48037));
    InMux I__11171 (
            .O(N__48042),
            .I(N__48037));
    LocalMux I__11170 (
            .O(N__48037),
            .I(N__48033));
    InMux I__11169 (
            .O(N__48036),
            .I(N__48030));
    Span4Mux_h I__11168 (
            .O(N__48033),
            .I(N__48027));
    LocalMux I__11167 (
            .O(N__48030),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__11166 (
            .O(N__48027),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__11165 (
            .O(N__48022),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__11164 (
            .O(N__48019),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__11163 (
            .O(N__48016),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__11162 (
            .O(N__48013),
            .I(N__48010));
    LocalMux I__11161 (
            .O(N__48010),
            .I(N__48006));
    InMux I__11160 (
            .O(N__48009),
            .I(N__48003));
    Span4Mux_v I__11159 (
            .O(N__48006),
            .I(N__48000));
    LocalMux I__11158 (
            .O(N__48003),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__11157 (
            .O(N__48000),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__11156 (
            .O(N__47995),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__11155 (
            .O(N__47992),
            .I(N__47989));
    LocalMux I__11154 (
            .O(N__47989),
            .I(N__47986));
    Span4Mux_v I__11153 (
            .O(N__47986),
            .I(N__47982));
    InMux I__11152 (
            .O(N__47985),
            .I(N__47979));
    Span4Mux_h I__11151 (
            .O(N__47982),
            .I(N__47976));
    LocalMux I__11150 (
            .O(N__47979),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__11149 (
            .O(N__47976),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__11148 (
            .O(N__47971),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__11147 (
            .O(N__47968),
            .I(N__47965));
    LocalMux I__11146 (
            .O(N__47965),
            .I(N__47962));
    Span4Mux_h I__11145 (
            .O(N__47962),
            .I(N__47958));
    InMux I__11144 (
            .O(N__47961),
            .I(N__47955));
    Span4Mux_v I__11143 (
            .O(N__47958),
            .I(N__47952));
    LocalMux I__11142 (
            .O(N__47955),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__11141 (
            .O(N__47952),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__11140 (
            .O(N__47947),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__11139 (
            .O(N__47944),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__11138 (
            .O(N__47941),
            .I(N__47937));
    InMux I__11137 (
            .O(N__47940),
            .I(N__47934));
    LocalMux I__11136 (
            .O(N__47937),
            .I(N__47931));
    LocalMux I__11135 (
            .O(N__47934),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv12 I__11134 (
            .O(N__47931),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__11133 (
            .O(N__47926),
            .I(bfn_18_14_0_));
    InMux I__11132 (
            .O(N__47923),
            .I(N__47919));
    InMux I__11131 (
            .O(N__47922),
            .I(N__47916));
    LocalMux I__11130 (
            .O(N__47919),
            .I(N__47913));
    LocalMux I__11129 (
            .O(N__47916),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv12 I__11128 (
            .O(N__47913),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__11127 (
            .O(N__47908),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__11126 (
            .O(N__47905),
            .I(N__47901));
    InMux I__11125 (
            .O(N__47904),
            .I(N__47898));
    LocalMux I__11124 (
            .O(N__47901),
            .I(N__47895));
    LocalMux I__11123 (
            .O(N__47898),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__11122 (
            .O(N__47895),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__11121 (
            .O(N__47890),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__11120 (
            .O(N__47887),
            .I(N__47883));
    InMux I__11119 (
            .O(N__47886),
            .I(N__47880));
    LocalMux I__11118 (
            .O(N__47883),
            .I(N__47877));
    LocalMux I__11117 (
            .O(N__47880),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__11116 (
            .O(N__47877),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__11115 (
            .O(N__47872),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__11114 (
            .O(N__47869),
            .I(N__47865));
    InMux I__11113 (
            .O(N__47868),
            .I(N__47862));
    LocalMux I__11112 (
            .O(N__47865),
            .I(N__47859));
    LocalMux I__11111 (
            .O(N__47862),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__11110 (
            .O(N__47859),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__11109 (
            .O(N__47854),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__11108 (
            .O(N__47851),
            .I(N__47847));
    InMux I__11107 (
            .O(N__47850),
            .I(N__47844));
    LocalMux I__11106 (
            .O(N__47847),
            .I(N__47841));
    LocalMux I__11105 (
            .O(N__47844),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__11104 (
            .O(N__47841),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__11103 (
            .O(N__47836),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__11102 (
            .O(N__47833),
            .I(N__47829));
    InMux I__11101 (
            .O(N__47832),
            .I(N__47826));
    LocalMux I__11100 (
            .O(N__47829),
            .I(N__47823));
    LocalMux I__11099 (
            .O(N__47826),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv12 I__11098 (
            .O(N__47823),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__11097 (
            .O(N__47818),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__11096 (
            .O(N__47815),
            .I(N__47808));
    InMux I__11095 (
            .O(N__47814),
            .I(N__47808));
    InMux I__11094 (
            .O(N__47813),
            .I(N__47805));
    LocalMux I__11093 (
            .O(N__47808),
            .I(N__47802));
    LocalMux I__11092 (
            .O(N__47805),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__11091 (
            .O(N__47802),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__11090 (
            .O(N__47797),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__11089 (
            .O(N__47794),
            .I(N__47786));
    InMux I__11088 (
            .O(N__47793),
            .I(N__47786));
    InMux I__11087 (
            .O(N__47792),
            .I(N__47781));
    InMux I__11086 (
            .O(N__47791),
            .I(N__47781));
    LocalMux I__11085 (
            .O(N__47786),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    LocalMux I__11084 (
            .O(N__47781),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ));
    CascadeMux I__11083 (
            .O(N__47776),
            .I(N__47772));
    InMux I__11082 (
            .O(N__47775),
            .I(N__47767));
    InMux I__11081 (
            .O(N__47772),
            .I(N__47767));
    LocalMux I__11080 (
            .O(N__47767),
            .I(N__47764));
    Span4Mux_h I__11079 (
            .O(N__47764),
            .I(N__47759));
    InMux I__11078 (
            .O(N__47763),
            .I(N__47756));
    InMux I__11077 (
            .O(N__47762),
            .I(N__47753));
    Odrv4 I__11076 (
            .O(N__47759),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    LocalMux I__11075 (
            .O(N__47756),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    LocalMux I__11074 (
            .O(N__47753),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ));
    CascadeMux I__11073 (
            .O(N__47746),
            .I(\delay_measurement_inst.delay_tr_timer.N_362_cascade_ ));
    InMux I__11072 (
            .O(N__47743),
            .I(N__47739));
    CascadeMux I__11071 (
            .O(N__47742),
            .I(N__47735));
    LocalMux I__11070 (
            .O(N__47739),
            .I(N__47731));
    InMux I__11069 (
            .O(N__47738),
            .I(N__47724));
    InMux I__11068 (
            .O(N__47735),
            .I(N__47724));
    InMux I__11067 (
            .O(N__47734),
            .I(N__47724));
    Odrv4 I__11066 (
            .O(N__47731),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    LocalMux I__11065 (
            .O(N__47724),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ));
    InMux I__11064 (
            .O(N__47719),
            .I(N__47715));
    InMux I__11063 (
            .O(N__47718),
            .I(N__47712));
    LocalMux I__11062 (
            .O(N__47715),
            .I(N__47708));
    LocalMux I__11061 (
            .O(N__47712),
            .I(N__47705));
    InMux I__11060 (
            .O(N__47711),
            .I(N__47702));
    Span4Mux_v I__11059 (
            .O(N__47708),
            .I(N__47697));
    Span4Mux_v I__11058 (
            .O(N__47705),
            .I(N__47697));
    LocalMux I__11057 (
            .O(N__47702),
            .I(N__47694));
    Odrv4 I__11056 (
            .O(N__47697),
            .I(\delay_measurement_inst.N_365 ));
    Odrv4 I__11055 (
            .O(N__47694),
            .I(\delay_measurement_inst.N_365 ));
    InMux I__11054 (
            .O(N__47689),
            .I(N__47686));
    LocalMux I__11053 (
            .O(N__47686),
            .I(N__47683));
    Odrv4 I__11052 (
            .O(N__47683),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    CascadeMux I__11051 (
            .O(N__47680),
            .I(N__47676));
    InMux I__11050 (
            .O(N__47679),
            .I(N__47673));
    InMux I__11049 (
            .O(N__47676),
            .I(N__47670));
    LocalMux I__11048 (
            .O(N__47673),
            .I(N__47664));
    LocalMux I__11047 (
            .O(N__47670),
            .I(N__47664));
    InMux I__11046 (
            .O(N__47669),
            .I(N__47661));
    Odrv4 I__11045 (
            .O(N__47664),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__11044 (
            .O(N__47661),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__11043 (
            .O(N__47656),
            .I(N__47652));
    InMux I__11042 (
            .O(N__47655),
            .I(N__47649));
    LocalMux I__11041 (
            .O(N__47652),
            .I(N__47646));
    LocalMux I__11040 (
            .O(N__47649),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv12 I__11039 (
            .O(N__47646),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__11038 (
            .O(N__47641),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__11037 (
            .O(N__47638),
            .I(N__47635));
    InMux I__11036 (
            .O(N__47635),
            .I(N__47632));
    LocalMux I__11035 (
            .O(N__47632),
            .I(N__47629));
    Span4Mux_h I__11034 (
            .O(N__47629),
            .I(N__47626));
    Odrv4 I__11033 (
            .O(N__47626),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28 ));
    InMux I__11032 (
            .O(N__47623),
            .I(N__47619));
    InMux I__11031 (
            .O(N__47622),
            .I(N__47616));
    LocalMux I__11030 (
            .O(N__47619),
            .I(N__47613));
    LocalMux I__11029 (
            .O(N__47616),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__11028 (
            .O(N__47613),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__11027 (
            .O(N__47608),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__11026 (
            .O(N__47605),
            .I(N__47602));
    LocalMux I__11025 (
            .O(N__47602),
            .I(N__47598));
    InMux I__11024 (
            .O(N__47601),
            .I(N__47595));
    Sp12to4 I__11023 (
            .O(N__47598),
            .I(N__47592));
    LocalMux I__11022 (
            .O(N__47595),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv12 I__11021 (
            .O(N__47592),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__11020 (
            .O(N__47587),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__11019 (
            .O(N__47584),
            .I(N__47580));
    InMux I__11018 (
            .O(N__47583),
            .I(N__47577));
    LocalMux I__11017 (
            .O(N__47580),
            .I(N__47574));
    LocalMux I__11016 (
            .O(N__47577),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv12 I__11015 (
            .O(N__47574),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__11014 (
            .O(N__47569),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__11013 (
            .O(N__47566),
            .I(N__47562));
    InMux I__11012 (
            .O(N__47565),
            .I(N__47559));
    LocalMux I__11011 (
            .O(N__47562),
            .I(N__47556));
    LocalMux I__11010 (
            .O(N__47559),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__11009 (
            .O(N__47556),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__11008 (
            .O(N__47551),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__11007 (
            .O(N__47548),
            .I(N__47545));
    LocalMux I__11006 (
            .O(N__47545),
            .I(N__47541));
    InMux I__11005 (
            .O(N__47544),
            .I(N__47538));
    Span4Mux_h I__11004 (
            .O(N__47541),
            .I(N__47535));
    LocalMux I__11003 (
            .O(N__47538),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__11002 (
            .O(N__47535),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__11001 (
            .O(N__47530),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__11000 (
            .O(N__47527),
            .I(N__47523));
    InMux I__10999 (
            .O(N__47526),
            .I(N__47520));
    LocalMux I__10998 (
            .O(N__47523),
            .I(N__47517));
    LocalMux I__10997 (
            .O(N__47520),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv12 I__10996 (
            .O(N__47517),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__10995 (
            .O(N__47512),
            .I(N__47508));
    InMux I__10994 (
            .O(N__47511),
            .I(N__47505));
    InMux I__10993 (
            .O(N__47508),
            .I(N__47502));
    LocalMux I__10992 (
            .O(N__47505),
            .I(N__47499));
    LocalMux I__10991 (
            .O(N__47502),
            .I(N__47495));
    Span4Mux_v I__10990 (
            .O(N__47499),
            .I(N__47492));
    InMux I__10989 (
            .O(N__47498),
            .I(N__47489));
    Span4Mux_v I__10988 (
            .O(N__47495),
            .I(N__47486));
    Odrv4 I__10987 (
            .O(N__47492),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__10986 (
            .O(N__47489),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv4 I__10985 (
            .O(N__47486),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    CEMux I__10984 (
            .O(N__47479),
            .I(N__47464));
    CEMux I__10983 (
            .O(N__47478),
            .I(N__47464));
    CEMux I__10982 (
            .O(N__47477),
            .I(N__47464));
    CEMux I__10981 (
            .O(N__47476),
            .I(N__47464));
    CEMux I__10980 (
            .O(N__47475),
            .I(N__47464));
    GlobalMux I__10979 (
            .O(N__47464),
            .I(N__47461));
    gio2CtrlBuf I__10978 (
            .O(N__47461),
            .I(\delay_measurement_inst.delay_tr_timer.N_399_i_g ));
    CascadeMux I__10977 (
            .O(N__47458),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ));
    CascadeMux I__10976 (
            .O(N__47455),
            .I(N__47452));
    InMux I__10975 (
            .O(N__47452),
            .I(N__47448));
    InMux I__10974 (
            .O(N__47451),
            .I(N__47445));
    LocalMux I__10973 (
            .O(N__47448),
            .I(N__47442));
    LocalMux I__10972 (
            .O(N__47445),
            .I(N__47439));
    Span4Mux_h I__10971 (
            .O(N__47442),
            .I(N__47436));
    Span4Mux_h I__10970 (
            .O(N__47439),
            .I(N__47433));
    Odrv4 I__10969 (
            .O(N__47436),
            .I(\delay_measurement_inst.delay_tr_timer.N_394 ));
    Odrv4 I__10968 (
            .O(N__47433),
            .I(\delay_measurement_inst.delay_tr_timer.N_394 ));
    InMux I__10967 (
            .O(N__47428),
            .I(N__47425));
    LocalMux I__10966 (
            .O(N__47425),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ));
    InMux I__10965 (
            .O(N__47422),
            .I(N__47418));
    InMux I__10964 (
            .O(N__47421),
            .I(N__47415));
    LocalMux I__10963 (
            .O(N__47418),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__10962 (
            .O(N__47415),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    CascadeMux I__10961 (
            .O(N__47410),
            .I(N__47407));
    InMux I__10960 (
            .O(N__47407),
            .I(N__47403));
    InMux I__10959 (
            .O(N__47406),
            .I(N__47400));
    LocalMux I__10958 (
            .O(N__47403),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__10957 (
            .O(N__47400),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__10956 (
            .O(N__47395),
            .I(N__47392));
    LocalMux I__10955 (
            .O(N__47392),
            .I(N__47389));
    Odrv4 I__10954 (
            .O(N__47389),
            .I(\delay_measurement_inst.delay_tr_timer.N_346 ));
    CascadeMux I__10953 (
            .O(N__47386),
            .I(N__47383));
    InMux I__10952 (
            .O(N__47383),
            .I(N__47378));
    InMux I__10951 (
            .O(N__47382),
            .I(N__47373));
    InMux I__10950 (
            .O(N__47381),
            .I(N__47373));
    LocalMux I__10949 (
            .O(N__47378),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__10948 (
            .O(N__47373),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    CascadeMux I__10947 (
            .O(N__47368),
            .I(N__47365));
    InMux I__10946 (
            .O(N__47365),
            .I(N__47361));
    CascadeMux I__10945 (
            .O(N__47364),
            .I(N__47358));
    LocalMux I__10944 (
            .O(N__47361),
            .I(N__47355));
    InMux I__10943 (
            .O(N__47358),
            .I(N__47352));
    Span12Mux_h I__10942 (
            .O(N__47355),
            .I(N__47348));
    LocalMux I__10941 (
            .O(N__47352),
            .I(N__47345));
    InMux I__10940 (
            .O(N__47351),
            .I(N__47342));
    Odrv12 I__10939 (
            .O(N__47348),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    Odrv4 I__10938 (
            .O(N__47345),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__10937 (
            .O(N__47342),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    CascadeMux I__10936 (
            .O(N__47335),
            .I(\delay_measurement_inst.delay_tr_timer.N_346_cascade_ ));
    CascadeMux I__10935 (
            .O(N__47332),
            .I(N__47329));
    InMux I__10934 (
            .O(N__47329),
            .I(N__47326));
    LocalMux I__10933 (
            .O(N__47326),
            .I(N__47323));
    Span4Mux_h I__10932 (
            .O(N__47323),
            .I(N__47319));
    InMux I__10931 (
            .O(N__47322),
            .I(N__47316));
    Odrv4 I__10930 (
            .O(N__47319),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__10929 (
            .O(N__47316),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__10928 (
            .O(N__47311),
            .I(N__47308));
    LocalMux I__10927 (
            .O(N__47308),
            .I(N__47305));
    Odrv4 I__10926 (
            .O(N__47305),
            .I(\delay_measurement_inst.delay_tr_timer.N_349 ));
    CascadeMux I__10925 (
            .O(N__47302),
            .I(N__47299));
    InMux I__10924 (
            .O(N__47299),
            .I(N__47296));
    LocalMux I__10923 (
            .O(N__47296),
            .I(N__47293));
    Span4Mux_h I__10922 (
            .O(N__47293),
            .I(N__47288));
    InMux I__10921 (
            .O(N__47292),
            .I(N__47285));
    InMux I__10920 (
            .O(N__47291),
            .I(N__47282));
    Odrv4 I__10919 (
            .O(N__47288),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__10918 (
            .O(N__47285),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    LocalMux I__10917 (
            .O(N__47282),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__10916 (
            .O(N__47275),
            .I(N__47272));
    LocalMux I__10915 (
            .O(N__47272),
            .I(N__47269));
    Span4Mux_h I__10914 (
            .O(N__47269),
            .I(N__47266));
    Span4Mux_h I__10913 (
            .O(N__47266),
            .I(N__47261));
    InMux I__10912 (
            .O(N__47265),
            .I(N__47258));
    InMux I__10911 (
            .O(N__47264),
            .I(N__47255));
    Odrv4 I__10910 (
            .O(N__47261),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    LocalMux I__10909 (
            .O(N__47258),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    LocalMux I__10908 (
            .O(N__47255),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    CascadeMux I__10907 (
            .O(N__47248),
            .I(\delay_measurement_inst.delay_tr_timer.N_349_cascade_ ));
    InMux I__10906 (
            .O(N__47245),
            .I(N__47242));
    LocalMux I__10905 (
            .O(N__47242),
            .I(N__47239));
    Span4Mux_h I__10904 (
            .O(N__47239),
            .I(N__47236));
    Odrv4 I__10903 (
            .O(N__47236),
            .I(\delay_measurement_inst.delay_tr_timer.N_351 ));
    InMux I__10902 (
            .O(N__47233),
            .I(N__47230));
    LocalMux I__10901 (
            .O(N__47230),
            .I(N__47227));
    Span4Mux_v I__10900 (
            .O(N__47227),
            .I(N__47222));
    InMux I__10899 (
            .O(N__47226),
            .I(N__47217));
    InMux I__10898 (
            .O(N__47225),
            .I(N__47217));
    Odrv4 I__10897 (
            .O(N__47222),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    LocalMux I__10896 (
            .O(N__47217),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__10895 (
            .O(N__47212),
            .I(N__47209));
    LocalMux I__10894 (
            .O(N__47209),
            .I(N__47204));
    InMux I__10893 (
            .O(N__47208),
            .I(N__47199));
    InMux I__10892 (
            .O(N__47207),
            .I(N__47199));
    Odrv4 I__10891 (
            .O(N__47204),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__10890 (
            .O(N__47199),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    CascadeMux I__10889 (
            .O(N__47194),
            .I(N__47190));
    InMux I__10888 (
            .O(N__47193),
            .I(N__47186));
    InMux I__10887 (
            .O(N__47190),
            .I(N__47183));
    InMux I__10886 (
            .O(N__47189),
            .I(N__47180));
    LocalMux I__10885 (
            .O(N__47186),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__10884 (
            .O(N__47183),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__10883 (
            .O(N__47180),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__10882 (
            .O(N__47173),
            .I(N__47168));
    InMux I__10881 (
            .O(N__47172),
            .I(N__47163));
    InMux I__10880 (
            .O(N__47171),
            .I(N__47163));
    LocalMux I__10879 (
            .O(N__47168),
            .I(N__47160));
    LocalMux I__10878 (
            .O(N__47163),
            .I(N__47157));
    Odrv12 I__10877 (
            .O(N__47160),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__10876 (
            .O(N__47157),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__10875 (
            .O(N__47152),
            .I(N__47149));
    LocalMux I__10874 (
            .O(N__47149),
            .I(N__47146));
    Span4Mux_h I__10873 (
            .O(N__47146),
            .I(N__47143));
    Odrv4 I__10872 (
            .O(N__47143),
            .I(\delay_measurement_inst.delay_tr_timer.N_362 ));
    InMux I__10871 (
            .O(N__47140),
            .I(N__47137));
    LocalMux I__10870 (
            .O(N__47137),
            .I(N__47134));
    Odrv12 I__10869 (
            .O(N__47134),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__10868 (
            .O(N__47131),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ));
    InMux I__10867 (
            .O(N__47128),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    InMux I__10866 (
            .O(N__47125),
            .I(N__47119));
    InMux I__10865 (
            .O(N__47124),
            .I(N__47119));
    LocalMux I__10864 (
            .O(N__47119),
            .I(N__47116));
    Odrv12 I__10863 (
            .O(N__47116),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__10862 (
            .O(N__47113),
            .I(N__47108));
    InMux I__10861 (
            .O(N__47112),
            .I(N__47102));
    InMux I__10860 (
            .O(N__47111),
            .I(N__47099));
    LocalMux I__10859 (
            .O(N__47108),
            .I(N__47094));
    InMux I__10858 (
            .O(N__47107),
            .I(N__47089));
    InMux I__10857 (
            .O(N__47106),
            .I(N__47089));
    CascadeMux I__10856 (
            .O(N__47105),
            .I(N__47080));
    LocalMux I__10855 (
            .O(N__47102),
            .I(N__47073));
    LocalMux I__10854 (
            .O(N__47099),
            .I(N__47052));
    InMux I__10853 (
            .O(N__47098),
            .I(N__47047));
    InMux I__10852 (
            .O(N__47097),
            .I(N__47047));
    Span4Mux_v I__10851 (
            .O(N__47094),
            .I(N__47042));
    LocalMux I__10850 (
            .O(N__47089),
            .I(N__47042));
    InMux I__10849 (
            .O(N__47088),
            .I(N__47033));
    InMux I__10848 (
            .O(N__47087),
            .I(N__47033));
    InMux I__10847 (
            .O(N__47086),
            .I(N__47033));
    InMux I__10846 (
            .O(N__47085),
            .I(N__47033));
    InMux I__10845 (
            .O(N__47084),
            .I(N__47028));
    InMux I__10844 (
            .O(N__47083),
            .I(N__47028));
    InMux I__10843 (
            .O(N__47080),
            .I(N__47021));
    InMux I__10842 (
            .O(N__47079),
            .I(N__47021));
    InMux I__10841 (
            .O(N__47078),
            .I(N__47021));
    InMux I__10840 (
            .O(N__47077),
            .I(N__47015));
    InMux I__10839 (
            .O(N__47076),
            .I(N__47015));
    Span4Mux_v I__10838 (
            .O(N__47073),
            .I(N__47012));
    InMux I__10837 (
            .O(N__47072),
            .I(N__46997));
    InMux I__10836 (
            .O(N__47071),
            .I(N__46997));
    InMux I__10835 (
            .O(N__47070),
            .I(N__46997));
    InMux I__10834 (
            .O(N__47069),
            .I(N__46997));
    InMux I__10833 (
            .O(N__47068),
            .I(N__46997));
    InMux I__10832 (
            .O(N__47067),
            .I(N__46997));
    InMux I__10831 (
            .O(N__47066),
            .I(N__46997));
    InMux I__10830 (
            .O(N__47065),
            .I(N__46986));
    InMux I__10829 (
            .O(N__47064),
            .I(N__46986));
    InMux I__10828 (
            .O(N__47063),
            .I(N__46986));
    InMux I__10827 (
            .O(N__47062),
            .I(N__46986));
    InMux I__10826 (
            .O(N__47061),
            .I(N__46986));
    InMux I__10825 (
            .O(N__47060),
            .I(N__46979));
    InMux I__10824 (
            .O(N__47059),
            .I(N__46979));
    InMux I__10823 (
            .O(N__47058),
            .I(N__46979));
    InMux I__10822 (
            .O(N__47057),
            .I(N__46972));
    InMux I__10821 (
            .O(N__47056),
            .I(N__46972));
    InMux I__10820 (
            .O(N__47055),
            .I(N__46972));
    Span4Mux_v I__10819 (
            .O(N__47052),
            .I(N__46959));
    LocalMux I__10818 (
            .O(N__47047),
            .I(N__46959));
    Span4Mux_h I__10817 (
            .O(N__47042),
            .I(N__46959));
    LocalMux I__10816 (
            .O(N__47033),
            .I(N__46959));
    LocalMux I__10815 (
            .O(N__47028),
            .I(N__46959));
    LocalMux I__10814 (
            .O(N__47021),
            .I(N__46959));
    InMux I__10813 (
            .O(N__47020),
            .I(N__46956));
    LocalMux I__10812 (
            .O(N__47015),
            .I(N__46951));
    Span4Mux_h I__10811 (
            .O(N__47012),
            .I(N__46951));
    LocalMux I__10810 (
            .O(N__46997),
            .I(N__46942));
    LocalMux I__10809 (
            .O(N__46986),
            .I(N__46942));
    LocalMux I__10808 (
            .O(N__46979),
            .I(N__46942));
    LocalMux I__10807 (
            .O(N__46972),
            .I(N__46942));
    Span4Mux_v I__10806 (
            .O(N__46959),
            .I(N__46939));
    LocalMux I__10805 (
            .O(N__46956),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    Odrv4 I__10804 (
            .O(N__46951),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    Odrv12 I__10803 (
            .O(N__46942),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    Odrv4 I__10802 (
            .O(N__46939),
            .I(elapsed_time_ns_1_RNI5IV8E1_0_31));
    CascadeMux I__10801 (
            .O(N__46930),
            .I(N__46919));
    InMux I__10800 (
            .O(N__46929),
            .I(N__46916));
    InMux I__10799 (
            .O(N__46928),
            .I(N__46905));
    InMux I__10798 (
            .O(N__46927),
            .I(N__46905));
    InMux I__10797 (
            .O(N__46926),
            .I(N__46905));
    InMux I__10796 (
            .O(N__46925),
            .I(N__46905));
    InMux I__10795 (
            .O(N__46924),
            .I(N__46905));
    InMux I__10794 (
            .O(N__46923),
            .I(N__46898));
    InMux I__10793 (
            .O(N__46922),
            .I(N__46898));
    InMux I__10792 (
            .O(N__46919),
            .I(N__46898));
    LocalMux I__10791 (
            .O(N__46916),
            .I(\phase_controller_inst1.stoper_hc.N_318 ));
    LocalMux I__10790 (
            .O(N__46905),
            .I(\phase_controller_inst1.stoper_hc.N_318 ));
    LocalMux I__10789 (
            .O(N__46898),
            .I(\phase_controller_inst1.stoper_hc.N_318 ));
    CascadeMux I__10788 (
            .O(N__46891),
            .I(N__46887));
    InMux I__10787 (
            .O(N__46890),
            .I(N__46881));
    InMux I__10786 (
            .O(N__46887),
            .I(N__46878));
    InMux I__10785 (
            .O(N__46886),
            .I(N__46875));
    InMux I__10784 (
            .O(N__46885),
            .I(N__46871));
    InMux I__10783 (
            .O(N__46884),
            .I(N__46867));
    LocalMux I__10782 (
            .O(N__46881),
            .I(N__46864));
    LocalMux I__10781 (
            .O(N__46878),
            .I(N__46861));
    LocalMux I__10780 (
            .O(N__46875),
            .I(N__46858));
    InMux I__10779 (
            .O(N__46874),
            .I(N__46855));
    LocalMux I__10778 (
            .O(N__46871),
            .I(N__46852));
    InMux I__10777 (
            .O(N__46870),
            .I(N__46849));
    LocalMux I__10776 (
            .O(N__46867),
            .I(N__46838));
    Span4Mux_v I__10775 (
            .O(N__46864),
            .I(N__46838));
    Span4Mux_v I__10774 (
            .O(N__46861),
            .I(N__46838));
    Span4Mux_v I__10773 (
            .O(N__46858),
            .I(N__46838));
    LocalMux I__10772 (
            .O(N__46855),
            .I(N__46838));
    Odrv4 I__10771 (
            .O(N__46852),
            .I(elapsed_time_ns_1_RNIDDC6P1_0_14));
    LocalMux I__10770 (
            .O(N__46849),
            .I(elapsed_time_ns_1_RNIDDC6P1_0_14));
    Odrv4 I__10769 (
            .O(N__46838),
            .I(elapsed_time_ns_1_RNIDDC6P1_0_14));
    CascadeMux I__10768 (
            .O(N__46831),
            .I(N__46819));
    CascadeMux I__10767 (
            .O(N__46830),
            .I(N__46816));
    CascadeMux I__10766 (
            .O(N__46829),
            .I(N__46813));
    InMux I__10765 (
            .O(N__46828),
            .I(N__46807));
    CascadeMux I__10764 (
            .O(N__46827),
            .I(N__46796));
    InMux I__10763 (
            .O(N__46826),
            .I(N__46791));
    InMux I__10762 (
            .O(N__46825),
            .I(N__46776));
    InMux I__10761 (
            .O(N__46824),
            .I(N__46776));
    InMux I__10760 (
            .O(N__46823),
            .I(N__46776));
    InMux I__10759 (
            .O(N__46822),
            .I(N__46776));
    InMux I__10758 (
            .O(N__46819),
            .I(N__46776));
    InMux I__10757 (
            .O(N__46816),
            .I(N__46776));
    InMux I__10756 (
            .O(N__46813),
            .I(N__46776));
    InMux I__10755 (
            .O(N__46812),
            .I(N__46773));
    InMux I__10754 (
            .O(N__46811),
            .I(N__46768));
    InMux I__10753 (
            .O(N__46810),
            .I(N__46768));
    LocalMux I__10752 (
            .O(N__46807),
            .I(N__46765));
    InMux I__10751 (
            .O(N__46806),
            .I(N__46754));
    InMux I__10750 (
            .O(N__46805),
            .I(N__46754));
    InMux I__10749 (
            .O(N__46804),
            .I(N__46754));
    InMux I__10748 (
            .O(N__46803),
            .I(N__46754));
    InMux I__10747 (
            .O(N__46802),
            .I(N__46754));
    InMux I__10746 (
            .O(N__46801),
            .I(N__46751));
    InMux I__10745 (
            .O(N__46800),
            .I(N__46748));
    InMux I__10744 (
            .O(N__46799),
            .I(N__46742));
    InMux I__10743 (
            .O(N__46796),
            .I(N__46735));
    InMux I__10742 (
            .O(N__46795),
            .I(N__46735));
    InMux I__10741 (
            .O(N__46794),
            .I(N__46735));
    LocalMux I__10740 (
            .O(N__46791),
            .I(N__46732));
    LocalMux I__10739 (
            .O(N__46776),
            .I(N__46729));
    LocalMux I__10738 (
            .O(N__46773),
            .I(N__46726));
    LocalMux I__10737 (
            .O(N__46768),
            .I(N__46719));
    Span4Mux_v I__10736 (
            .O(N__46765),
            .I(N__46719));
    LocalMux I__10735 (
            .O(N__46754),
            .I(N__46719));
    LocalMux I__10734 (
            .O(N__46751),
            .I(N__46714));
    LocalMux I__10733 (
            .O(N__46748),
            .I(N__46714));
    InMux I__10732 (
            .O(N__46747),
            .I(N__46709));
    InMux I__10731 (
            .O(N__46746),
            .I(N__46709));
    InMux I__10730 (
            .O(N__46745),
            .I(N__46706));
    LocalMux I__10729 (
            .O(N__46742),
            .I(N__46699));
    LocalMux I__10728 (
            .O(N__46735),
            .I(N__46699));
    Span4Mux_h I__10727 (
            .O(N__46732),
            .I(N__46699));
    Span4Mux_v I__10726 (
            .O(N__46729),
            .I(N__46694));
    Span4Mux_h I__10725 (
            .O(N__46726),
            .I(N__46694));
    Span4Mux_v I__10724 (
            .O(N__46719),
            .I(N__46687));
    Span4Mux_v I__10723 (
            .O(N__46714),
            .I(N__46687));
    LocalMux I__10722 (
            .O(N__46709),
            .I(N__46687));
    LocalMux I__10721 (
            .O(N__46706),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    Odrv4 I__10720 (
            .O(N__46699),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    Odrv4 I__10719 (
            .O(N__46694),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    Odrv4 I__10718 (
            .O(N__46687),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ));
    CascadeMux I__10717 (
            .O(N__46678),
            .I(N__46675));
    InMux I__10716 (
            .O(N__46675),
            .I(N__46672));
    LocalMux I__10715 (
            .O(N__46672),
            .I(N__46669));
    Odrv12 I__10714 (
            .O(N__46669),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    InMux I__10713 (
            .O(N__46666),
            .I(N__46660));
    InMux I__10712 (
            .O(N__46665),
            .I(N__46657));
    InMux I__10711 (
            .O(N__46664),
            .I(N__46653));
    InMux I__10710 (
            .O(N__46663),
            .I(N__46650));
    LocalMux I__10709 (
            .O(N__46660),
            .I(N__46647));
    LocalMux I__10708 (
            .O(N__46657),
            .I(N__46644));
    CascadeMux I__10707 (
            .O(N__46656),
            .I(N__46640));
    LocalMux I__10706 (
            .O(N__46653),
            .I(N__46635));
    LocalMux I__10705 (
            .O(N__46650),
            .I(N__46635));
    Span4Mux_v I__10704 (
            .O(N__46647),
            .I(N__46632));
    Sp12to4 I__10703 (
            .O(N__46644),
            .I(N__46629));
    InMux I__10702 (
            .O(N__46643),
            .I(N__46626));
    InMux I__10701 (
            .O(N__46640),
            .I(N__46623));
    Span4Mux_v I__10700 (
            .O(N__46635),
            .I(N__46618));
    Span4Mux_h I__10699 (
            .O(N__46632),
            .I(N__46618));
    Span12Mux_h I__10698 (
            .O(N__46629),
            .I(N__46615));
    LocalMux I__10697 (
            .O(N__46626),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__10696 (
            .O(N__46623),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__10695 (
            .O(N__46618),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__10694 (
            .O(N__46615),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    CascadeMux I__10693 (
            .O(N__46606),
            .I(N__46603));
    InMux I__10692 (
            .O(N__46603),
            .I(N__46600));
    LocalMux I__10691 (
            .O(N__46600),
            .I(N__46595));
    InMux I__10690 (
            .O(N__46599),
            .I(N__46592));
    InMux I__10689 (
            .O(N__46598),
            .I(N__46589));
    Span4Mux_h I__10688 (
            .O(N__46595),
            .I(N__46584));
    LocalMux I__10687 (
            .O(N__46592),
            .I(N__46581));
    LocalMux I__10686 (
            .O(N__46589),
            .I(N__46578));
    InMux I__10685 (
            .O(N__46588),
            .I(N__46575));
    InMux I__10684 (
            .O(N__46587),
            .I(N__46572));
    Span4Mux_v I__10683 (
            .O(N__46584),
            .I(N__46569));
    Span4Mux_h I__10682 (
            .O(N__46581),
            .I(N__46564));
    Span4Mux_h I__10681 (
            .O(N__46578),
            .I(N__46564));
    LocalMux I__10680 (
            .O(N__46575),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__10679 (
            .O(N__46572),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__10678 (
            .O(N__46569),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__10677 (
            .O(N__46564),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    IoInMux I__10676 (
            .O(N__46555),
            .I(N__46552));
    LocalMux I__10675 (
            .O(N__46552),
            .I(N__46549));
    Span4Mux_s1_v I__10674 (
            .O(N__46549),
            .I(N__46546));
    Span4Mux_v I__10673 (
            .O(N__46546),
            .I(N__46542));
    InMux I__10672 (
            .O(N__46545),
            .I(N__46539));
    Odrv4 I__10671 (
            .O(N__46542),
            .I(T12_c));
    LocalMux I__10670 (
            .O(N__46539),
            .I(T12_c));
    CascadeMux I__10669 (
            .O(N__46534),
            .I(N__46530));
    InMux I__10668 (
            .O(N__46533),
            .I(N__46527));
    InMux I__10667 (
            .O(N__46530),
            .I(N__46524));
    LocalMux I__10666 (
            .O(N__46527),
            .I(N__46521));
    LocalMux I__10665 (
            .O(N__46524),
            .I(N__46517));
    Span4Mux_v I__10664 (
            .O(N__46521),
            .I(N__46514));
    InMux I__10663 (
            .O(N__46520),
            .I(N__46511));
    Span4Mux_v I__10662 (
            .O(N__46517),
            .I(N__46508));
    Odrv4 I__10661 (
            .O(N__46514),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__10660 (
            .O(N__46511),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__10659 (
            .O(N__46508),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    CascadeMux I__10658 (
            .O(N__46501),
            .I(N__46498));
    InMux I__10657 (
            .O(N__46498),
            .I(N__46495));
    LocalMux I__10656 (
            .O(N__46495),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__10655 (
            .O(N__46492),
            .I(N__46489));
    LocalMux I__10654 (
            .O(N__46489),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__10653 (
            .O(N__46486),
            .I(N__46483));
    LocalMux I__10652 (
            .O(N__46483),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    CascadeMux I__10651 (
            .O(N__46480),
            .I(N__46477));
    InMux I__10650 (
            .O(N__46477),
            .I(N__46474));
    LocalMux I__10649 (
            .O(N__46474),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__10648 (
            .O(N__46471),
            .I(N__46468));
    LocalMux I__10647 (
            .O(N__46468),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__10646 (
            .O(N__46465),
            .I(N__46462));
    LocalMux I__10645 (
            .O(N__46462),
            .I(N__46459));
    Odrv4 I__10644 (
            .O(N__46459),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__10643 (
            .O(N__46456),
            .I(N__46453));
    InMux I__10642 (
            .O(N__46453),
            .I(N__46450));
    LocalMux I__10641 (
            .O(N__46450),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__10640 (
            .O(N__46447),
            .I(N__46444));
    LocalMux I__10639 (
            .O(N__46444),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    CascadeMux I__10638 (
            .O(N__46441),
            .I(N__46438));
    InMux I__10637 (
            .O(N__46438),
            .I(N__46435));
    LocalMux I__10636 (
            .O(N__46435),
            .I(N__46432));
    Odrv4 I__10635 (
            .O(N__46432),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    InMux I__10634 (
            .O(N__46429),
            .I(N__46426));
    LocalMux I__10633 (
            .O(N__46426),
            .I(N__46423));
    Odrv4 I__10632 (
            .O(N__46423),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    CascadeMux I__10631 (
            .O(N__46420),
            .I(N__46417));
    InMux I__10630 (
            .O(N__46417),
            .I(N__46414));
    LocalMux I__10629 (
            .O(N__46414),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    InMux I__10628 (
            .O(N__46411),
            .I(N__46408));
    LocalMux I__10627 (
            .O(N__46408),
            .I(N__46405));
    Odrv12 I__10626 (
            .O(N__46405),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__10625 (
            .O(N__46402),
            .I(N__46399));
    InMux I__10624 (
            .O(N__46399),
            .I(N__46396));
    LocalMux I__10623 (
            .O(N__46396),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__10622 (
            .O(N__46393),
            .I(N__46390));
    LocalMux I__10621 (
            .O(N__46390),
            .I(N__46387));
    Span4Mux_v I__10620 (
            .O(N__46387),
            .I(N__46384));
    Odrv4 I__10619 (
            .O(N__46384),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__10618 (
            .O(N__46381),
            .I(N__46378));
    InMux I__10617 (
            .O(N__46378),
            .I(N__46375));
    LocalMux I__10616 (
            .O(N__46375),
            .I(N__46372));
    Odrv4 I__10615 (
            .O(N__46372),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__10614 (
            .O(N__46369),
            .I(N__46366));
    LocalMux I__10613 (
            .O(N__46366),
            .I(N__46363));
    Span4Mux_v I__10612 (
            .O(N__46363),
            .I(N__46360));
    Span4Mux_h I__10611 (
            .O(N__46360),
            .I(N__46357));
    Odrv4 I__10610 (
            .O(N__46357),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__10609 (
            .O(N__46354),
            .I(N__46351));
    InMux I__10608 (
            .O(N__46351),
            .I(N__46348));
    LocalMux I__10607 (
            .O(N__46348),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    InMux I__10606 (
            .O(N__46345),
            .I(N__46342));
    LocalMux I__10605 (
            .O(N__46342),
            .I(N__46339));
    Span4Mux_v I__10604 (
            .O(N__46339),
            .I(N__46336));
    Span4Mux_h I__10603 (
            .O(N__46336),
            .I(N__46333));
    Odrv4 I__10602 (
            .O(N__46333),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    CascadeMux I__10601 (
            .O(N__46330),
            .I(N__46327));
    InMux I__10600 (
            .O(N__46327),
            .I(N__46324));
    LocalMux I__10599 (
            .O(N__46324),
            .I(N__46321));
    Odrv4 I__10598 (
            .O(N__46321),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__10597 (
            .O(N__46318),
            .I(N__46315));
    LocalMux I__10596 (
            .O(N__46315),
            .I(N__46312));
    Odrv12 I__10595 (
            .O(N__46312),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__10594 (
            .O(N__46309),
            .I(N__46306));
    InMux I__10593 (
            .O(N__46306),
            .I(N__46303));
    LocalMux I__10592 (
            .O(N__46303),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__10591 (
            .O(N__46300),
            .I(N__46297));
    LocalMux I__10590 (
            .O(N__46297),
            .I(N__46294));
    Odrv4 I__10589 (
            .O(N__46294),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__10588 (
            .O(N__46291),
            .I(N__46288));
    InMux I__10587 (
            .O(N__46288),
            .I(N__46285));
    LocalMux I__10586 (
            .O(N__46285),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__10585 (
            .O(N__46282),
            .I(N__46279));
    LocalMux I__10584 (
            .O(N__46279),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__10583 (
            .O(N__46276),
            .I(N__46273));
    InMux I__10582 (
            .O(N__46273),
            .I(N__46270));
    LocalMux I__10581 (
            .O(N__46270),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__10580 (
            .O(N__46267),
            .I(N__46264));
    LocalMux I__10579 (
            .O(N__46264),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__10578 (
            .O(N__46261),
            .I(N__46258));
    InMux I__10577 (
            .O(N__46258),
            .I(N__46255));
    LocalMux I__10576 (
            .O(N__46255),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__10575 (
            .O(N__46252),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__10574 (
            .O(N__46249),
            .I(N__46246));
    InMux I__10573 (
            .O(N__46246),
            .I(N__46240));
    InMux I__10572 (
            .O(N__46245),
            .I(N__46240));
    LocalMux I__10571 (
            .O(N__46240),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__10570 (
            .O(N__46237),
            .I(N__46234));
    InMux I__10569 (
            .O(N__46234),
            .I(N__46228));
    InMux I__10568 (
            .O(N__46233),
            .I(N__46228));
    LocalMux I__10567 (
            .O(N__46228),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    CascadeMux I__10566 (
            .O(N__46225),
            .I(N__46222));
    InMux I__10565 (
            .O(N__46222),
            .I(N__46215));
    InMux I__10564 (
            .O(N__46221),
            .I(N__46206));
    InMux I__10563 (
            .O(N__46220),
            .I(N__46206));
    InMux I__10562 (
            .O(N__46219),
            .I(N__46206));
    InMux I__10561 (
            .O(N__46218),
            .I(N__46206));
    LocalMux I__10560 (
            .O(N__46215),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    LocalMux I__10559 (
            .O(N__46206),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    CascadeMux I__10558 (
            .O(N__46201),
            .I(N__46198));
    InMux I__10557 (
            .O(N__46198),
            .I(N__46194));
    CascadeMux I__10556 (
            .O(N__46197),
            .I(N__46191));
    LocalMux I__10555 (
            .O(N__46194),
            .I(N__46187));
    InMux I__10554 (
            .O(N__46191),
            .I(N__46182));
    InMux I__10553 (
            .O(N__46190),
            .I(N__46182));
    Span4Mux_v I__10552 (
            .O(N__46187),
            .I(N__46178));
    LocalMux I__10551 (
            .O(N__46182),
            .I(N__46175));
    InMux I__10550 (
            .O(N__46181),
            .I(N__46172));
    Span4Mux_h I__10549 (
            .O(N__46178),
            .I(N__46169));
    Span4Mux_v I__10548 (
            .O(N__46175),
            .I(N__46166));
    LocalMux I__10547 (
            .O(N__46172),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__10546 (
            .O(N__46169),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv4 I__10545 (
            .O(N__46166),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__10544 (
            .O(N__46159),
            .I(N__46153));
    InMux I__10543 (
            .O(N__46158),
            .I(N__46153));
    LocalMux I__10542 (
            .O(N__46153),
            .I(N__46148));
    InMux I__10541 (
            .O(N__46152),
            .I(N__46143));
    InMux I__10540 (
            .O(N__46151),
            .I(N__46143));
    Span4Mux_v I__10539 (
            .O(N__46148),
            .I(N__46140));
    LocalMux I__10538 (
            .O(N__46143),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__10537 (
            .O(N__46140),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__10536 (
            .O(N__46135),
            .I(N__46132));
    LocalMux I__10535 (
            .O(N__46132),
            .I(N__46129));
    Span4Mux_v I__10534 (
            .O(N__46129),
            .I(N__46122));
    InMux I__10533 (
            .O(N__46128),
            .I(N__46113));
    InMux I__10532 (
            .O(N__46127),
            .I(N__46113));
    InMux I__10531 (
            .O(N__46126),
            .I(N__46113));
    InMux I__10530 (
            .O(N__46125),
            .I(N__46113));
    Odrv4 I__10529 (
            .O(N__46122),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__10528 (
            .O(N__46113),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    InMux I__10527 (
            .O(N__46108),
            .I(N__46105));
    LocalMux I__10526 (
            .O(N__46105),
            .I(N__46102));
    Odrv12 I__10525 (
            .O(N__46102),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__10524 (
            .O(N__46099),
            .I(N__46096));
    InMux I__10523 (
            .O(N__46096),
            .I(N__46093));
    LocalMux I__10522 (
            .O(N__46093),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__10521 (
            .O(N__46090),
            .I(N__46087));
    LocalMux I__10520 (
            .O(N__46087),
            .I(N__46084));
    Span4Mux_h I__10519 (
            .O(N__46084),
            .I(N__46081));
    Odrv4 I__10518 (
            .O(N__46081),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__10517 (
            .O(N__46078),
            .I(N__46075));
    InMux I__10516 (
            .O(N__46075),
            .I(N__46072));
    LocalMux I__10515 (
            .O(N__46072),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    InMux I__10514 (
            .O(N__46069),
            .I(N__46066));
    LocalMux I__10513 (
            .O(N__46066),
            .I(N__46063));
    Span4Mux_h I__10512 (
            .O(N__46063),
            .I(N__46060));
    Odrv4 I__10511 (
            .O(N__46060),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__10510 (
            .O(N__46057),
            .I(N__46054));
    InMux I__10509 (
            .O(N__46054),
            .I(N__46051));
    LocalMux I__10508 (
            .O(N__46051),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__10507 (
            .O(N__46048),
            .I(N__46044));
    InMux I__10506 (
            .O(N__46047),
            .I(N__46041));
    LocalMux I__10505 (
            .O(N__46044),
            .I(N__46038));
    LocalMux I__10504 (
            .O(N__46041),
            .I(N__46035));
    Span4Mux_h I__10503 (
            .O(N__46038),
            .I(N__46032));
    Odrv4 I__10502 (
            .O(N__46035),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    Odrv4 I__10501 (
            .O(N__46032),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    CascadeMux I__10500 (
            .O(N__46027),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_ ));
    InMux I__10499 (
            .O(N__46024),
            .I(N__46020));
    InMux I__10498 (
            .O(N__46023),
            .I(N__46017));
    LocalMux I__10497 (
            .O(N__46020),
            .I(N__46008));
    LocalMux I__10496 (
            .O(N__46017),
            .I(N__46008));
    InMux I__10495 (
            .O(N__46016),
            .I(N__46005));
    InMux I__10494 (
            .O(N__46015),
            .I(N__46001));
    InMux I__10493 (
            .O(N__46014),
            .I(N__45997));
    InMux I__10492 (
            .O(N__46013),
            .I(N__45994));
    Span4Mux_h I__10491 (
            .O(N__46008),
            .I(N__45991));
    LocalMux I__10490 (
            .O(N__46005),
            .I(N__45988));
    InMux I__10489 (
            .O(N__46004),
            .I(N__45985));
    LocalMux I__10488 (
            .O(N__46001),
            .I(N__45982));
    InMux I__10487 (
            .O(N__46000),
            .I(N__45979));
    LocalMux I__10486 (
            .O(N__45997),
            .I(\delay_measurement_inst.delay_hc_timer.N_344_i ));
    LocalMux I__10485 (
            .O(N__45994),
            .I(\delay_measurement_inst.delay_hc_timer.N_344_i ));
    Odrv4 I__10484 (
            .O(N__45991),
            .I(\delay_measurement_inst.delay_hc_timer.N_344_i ));
    Odrv4 I__10483 (
            .O(N__45988),
            .I(\delay_measurement_inst.delay_hc_timer.N_344_i ));
    LocalMux I__10482 (
            .O(N__45985),
            .I(\delay_measurement_inst.delay_hc_timer.N_344_i ));
    Odrv12 I__10481 (
            .O(N__45982),
            .I(\delay_measurement_inst.delay_hc_timer.N_344_i ));
    LocalMux I__10480 (
            .O(N__45979),
            .I(\delay_measurement_inst.delay_hc_timer.N_344_i ));
    InMux I__10479 (
            .O(N__45964),
            .I(N__45961));
    LocalMux I__10478 (
            .O(N__45961),
            .I(N__45955));
    InMux I__10477 (
            .O(N__45960),
            .I(N__45950));
    InMux I__10476 (
            .O(N__45959),
            .I(N__45950));
    InMux I__10475 (
            .O(N__45958),
            .I(N__45947));
    Span12Mux_v I__10474 (
            .O(N__45955),
            .I(N__45942));
    LocalMux I__10473 (
            .O(N__45950),
            .I(N__45942));
    LocalMux I__10472 (
            .O(N__45947),
            .I(elapsed_time_ns_1_RNIUE3CP1_0_6));
    Odrv12 I__10471 (
            .O(N__45942),
            .I(elapsed_time_ns_1_RNIUE3CP1_0_6));
    InMux I__10470 (
            .O(N__45937),
            .I(N__45933));
    CascadeMux I__10469 (
            .O(N__45936),
            .I(N__45930));
    LocalMux I__10468 (
            .O(N__45933),
            .I(N__45923));
    InMux I__10467 (
            .O(N__45930),
            .I(N__45919));
    InMux I__10466 (
            .O(N__45929),
            .I(N__45916));
    CascadeMux I__10465 (
            .O(N__45928),
            .I(N__45912));
    CascadeMux I__10464 (
            .O(N__45927),
            .I(N__45908));
    InMux I__10463 (
            .O(N__45926),
            .I(N__45899));
    Span4Mux_v I__10462 (
            .O(N__45923),
            .I(N__45896));
    InMux I__10461 (
            .O(N__45922),
            .I(N__45893));
    LocalMux I__10460 (
            .O(N__45919),
            .I(N__45888));
    LocalMux I__10459 (
            .O(N__45916),
            .I(N__45888));
    InMux I__10458 (
            .O(N__45915),
            .I(N__45881));
    InMux I__10457 (
            .O(N__45912),
            .I(N__45881));
    InMux I__10456 (
            .O(N__45911),
            .I(N__45881));
    InMux I__10455 (
            .O(N__45908),
            .I(N__45878));
    CascadeMux I__10454 (
            .O(N__45907),
            .I(N__45875));
    CascadeMux I__10453 (
            .O(N__45906),
            .I(N__45869));
    CascadeMux I__10452 (
            .O(N__45905),
            .I(N__45865));
    CascadeMux I__10451 (
            .O(N__45904),
            .I(N__45862));
    InMux I__10450 (
            .O(N__45903),
            .I(N__45855));
    InMux I__10449 (
            .O(N__45902),
            .I(N__45855));
    LocalMux I__10448 (
            .O(N__45899),
            .I(N__45848));
    Span4Mux_h I__10447 (
            .O(N__45896),
            .I(N__45848));
    LocalMux I__10446 (
            .O(N__45893),
            .I(N__45848));
    Span4Mux_h I__10445 (
            .O(N__45888),
            .I(N__45841));
    LocalMux I__10444 (
            .O(N__45881),
            .I(N__45841));
    LocalMux I__10443 (
            .O(N__45878),
            .I(N__45841));
    InMux I__10442 (
            .O(N__45875),
            .I(N__45830));
    InMux I__10441 (
            .O(N__45874),
            .I(N__45830));
    InMux I__10440 (
            .O(N__45873),
            .I(N__45830));
    InMux I__10439 (
            .O(N__45872),
            .I(N__45830));
    InMux I__10438 (
            .O(N__45869),
            .I(N__45830));
    InMux I__10437 (
            .O(N__45868),
            .I(N__45819));
    InMux I__10436 (
            .O(N__45865),
            .I(N__45819));
    InMux I__10435 (
            .O(N__45862),
            .I(N__45819));
    InMux I__10434 (
            .O(N__45861),
            .I(N__45819));
    InMux I__10433 (
            .O(N__45860),
            .I(N__45819));
    LocalMux I__10432 (
            .O(N__45855),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    Odrv4 I__10431 (
            .O(N__45848),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    Odrv4 I__10430 (
            .O(N__45841),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    LocalMux I__10429 (
            .O(N__45830),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    LocalMux I__10428 (
            .O(N__45819),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ));
    InMux I__10427 (
            .O(N__45808),
            .I(N__45805));
    LocalMux I__10426 (
            .O(N__45805),
            .I(N__45802));
    Span4Mux_h I__10425 (
            .O(N__45802),
            .I(N__45798));
    InMux I__10424 (
            .O(N__45801),
            .I(N__45795));
    Odrv4 I__10423 (
            .O(N__45798),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    LocalMux I__10422 (
            .O(N__45795),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    CascadeMux I__10421 (
            .O(N__45790),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15_cascade_));
    InMux I__10420 (
            .O(N__45787),
            .I(N__45783));
    InMux I__10419 (
            .O(N__45786),
            .I(N__45780));
    LocalMux I__10418 (
            .O(N__45783),
            .I(N__45774));
    LocalMux I__10417 (
            .O(N__45780),
            .I(N__45774));
    InMux I__10416 (
            .O(N__45779),
            .I(N__45771));
    Span4Mux_v I__10415 (
            .O(N__45774),
            .I(N__45768));
    LocalMux I__10414 (
            .O(N__45771),
            .I(N__45765));
    Span4Mux_h I__10413 (
            .O(N__45768),
            .I(N__45762));
    Odrv4 I__10412 (
            .O(N__45765),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ));
    Odrv4 I__10411 (
            .O(N__45762),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ));
    InMux I__10410 (
            .O(N__45757),
            .I(N__45753));
    InMux I__10409 (
            .O(N__45756),
            .I(N__45750));
    LocalMux I__10408 (
            .O(N__45753),
            .I(N__45747));
    LocalMux I__10407 (
            .O(N__45750),
            .I(N__45744));
    Span4Mux_h I__10406 (
            .O(N__45747),
            .I(N__45739));
    Span4Mux_v I__10405 (
            .O(N__45744),
            .I(N__45739));
    Odrv4 I__10404 (
            .O(N__45739),
            .I(\phase_controller_inst1.stoper_hc.N_269_iZ0Z_1 ));
    CascadeMux I__10403 (
            .O(N__45736),
            .I(N__45732));
    InMux I__10402 (
            .O(N__45735),
            .I(N__45727));
    InMux I__10401 (
            .O(N__45732),
            .I(N__45724));
    InMux I__10400 (
            .O(N__45731),
            .I(N__45721));
    CascadeMux I__10399 (
            .O(N__45730),
            .I(N__45718));
    LocalMux I__10398 (
            .O(N__45727),
            .I(N__45714));
    LocalMux I__10397 (
            .O(N__45724),
            .I(N__45709));
    LocalMux I__10396 (
            .O(N__45721),
            .I(N__45709));
    InMux I__10395 (
            .O(N__45718),
            .I(N__45706));
    CascadeMux I__10394 (
            .O(N__45717),
            .I(N__45702));
    Span4Mux_v I__10393 (
            .O(N__45714),
            .I(N__45694));
    Span4Mux_v I__10392 (
            .O(N__45709),
            .I(N__45694));
    LocalMux I__10391 (
            .O(N__45706),
            .I(N__45694));
    InMux I__10390 (
            .O(N__45705),
            .I(N__45691));
    InMux I__10389 (
            .O(N__45702),
            .I(N__45686));
    InMux I__10388 (
            .O(N__45701),
            .I(N__45686));
    Span4Mux_h I__10387 (
            .O(N__45694),
            .I(N__45683));
    LocalMux I__10386 (
            .O(N__45691),
            .I(N__45680));
    LocalMux I__10385 (
            .O(N__45686),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15));
    Odrv4 I__10384 (
            .O(N__45683),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15));
    Odrv12 I__10383 (
            .O(N__45680),
            .I(elapsed_time_ns_1_RNI7IT8E1_0_15));
    InMux I__10382 (
            .O(N__45673),
            .I(N__45669));
    InMux I__10381 (
            .O(N__45672),
            .I(N__45665));
    LocalMux I__10380 (
            .O(N__45669),
            .I(N__45662));
    InMux I__10379 (
            .O(N__45668),
            .I(N__45659));
    LocalMux I__10378 (
            .O(N__45665),
            .I(N__45656));
    Span4Mux_v I__10377 (
            .O(N__45662),
            .I(N__45649));
    LocalMux I__10376 (
            .O(N__45659),
            .I(N__45649));
    Span4Mux_h I__10375 (
            .O(N__45656),
            .I(N__45646));
    InMux I__10374 (
            .O(N__45655),
            .I(N__45641));
    InMux I__10373 (
            .O(N__45654),
            .I(N__45641));
    Span4Mux_h I__10372 (
            .O(N__45649),
            .I(N__45638));
    Odrv4 I__10371 (
            .O(N__45646),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    LocalMux I__10370 (
            .O(N__45641),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    Odrv4 I__10369 (
            .O(N__45638),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ));
    CascadeMux I__10368 (
            .O(N__45631),
            .I(N__45627));
    InMux I__10367 (
            .O(N__45630),
            .I(N__45624));
    InMux I__10366 (
            .O(N__45627),
            .I(N__45621));
    LocalMux I__10365 (
            .O(N__45624),
            .I(N__45618));
    LocalMux I__10364 (
            .O(N__45621),
            .I(N__45615));
    Odrv4 I__10363 (
            .O(N__45618),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv12 I__10362 (
            .O(N__45615),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    CascadeMux I__10361 (
            .O(N__45610),
            .I(N__45606));
    InMux I__10360 (
            .O(N__45609),
            .I(N__45603));
    InMux I__10359 (
            .O(N__45606),
            .I(N__45599));
    LocalMux I__10358 (
            .O(N__45603),
            .I(N__45596));
    CascadeMux I__10357 (
            .O(N__45602),
            .I(N__45593));
    LocalMux I__10356 (
            .O(N__45599),
            .I(N__45590));
    Span4Mux_v I__10355 (
            .O(N__45596),
            .I(N__45585));
    InMux I__10354 (
            .O(N__45593),
            .I(N__45582));
    Span4Mux_h I__10353 (
            .O(N__45590),
            .I(N__45579));
    InMux I__10352 (
            .O(N__45589),
            .I(N__45576));
    InMux I__10351 (
            .O(N__45588),
            .I(N__45573));
    Odrv4 I__10350 (
            .O(N__45585),
            .I(elapsed_time_ns_1_RNI1I3CP1_0_9));
    LocalMux I__10349 (
            .O(N__45582),
            .I(elapsed_time_ns_1_RNI1I3CP1_0_9));
    Odrv4 I__10348 (
            .O(N__45579),
            .I(elapsed_time_ns_1_RNI1I3CP1_0_9));
    LocalMux I__10347 (
            .O(N__45576),
            .I(elapsed_time_ns_1_RNI1I3CP1_0_9));
    LocalMux I__10346 (
            .O(N__45573),
            .I(elapsed_time_ns_1_RNI1I3CP1_0_9));
    CascadeMux I__10345 (
            .O(N__45562),
            .I(N__45557));
    InMux I__10344 (
            .O(N__45561),
            .I(N__45553));
    InMux I__10343 (
            .O(N__45560),
            .I(N__45540));
    InMux I__10342 (
            .O(N__45557),
            .I(N__45540));
    CascadeMux I__10341 (
            .O(N__45556),
            .I(N__45537));
    LocalMux I__10340 (
            .O(N__45553),
            .I(N__45534));
    CascadeMux I__10339 (
            .O(N__45552),
            .I(N__45531));
    CascadeMux I__10338 (
            .O(N__45551),
            .I(N__45528));
    CascadeMux I__10337 (
            .O(N__45550),
            .I(N__45525));
    CascadeMux I__10336 (
            .O(N__45549),
            .I(N__45521));
    InMux I__10335 (
            .O(N__45548),
            .I(N__45518));
    InMux I__10334 (
            .O(N__45547),
            .I(N__45515));
    InMux I__10333 (
            .O(N__45546),
            .I(N__45508));
    InMux I__10332 (
            .O(N__45545),
            .I(N__45505));
    LocalMux I__10331 (
            .O(N__45540),
            .I(N__45502));
    InMux I__10330 (
            .O(N__45537),
            .I(N__45499));
    Span4Mux_v I__10329 (
            .O(N__45534),
            .I(N__45496));
    InMux I__10328 (
            .O(N__45531),
            .I(N__45491));
    InMux I__10327 (
            .O(N__45528),
            .I(N__45491));
    InMux I__10326 (
            .O(N__45525),
            .I(N__45486));
    InMux I__10325 (
            .O(N__45524),
            .I(N__45486));
    InMux I__10324 (
            .O(N__45521),
            .I(N__45483));
    LocalMux I__10323 (
            .O(N__45518),
            .I(N__45478));
    LocalMux I__10322 (
            .O(N__45515),
            .I(N__45478));
    InMux I__10321 (
            .O(N__45514),
            .I(N__45471));
    InMux I__10320 (
            .O(N__45513),
            .I(N__45471));
    InMux I__10319 (
            .O(N__45512),
            .I(N__45471));
    CascadeMux I__10318 (
            .O(N__45511),
            .I(N__45467));
    LocalMux I__10317 (
            .O(N__45508),
            .I(N__45450));
    LocalMux I__10316 (
            .O(N__45505),
            .I(N__45450));
    Span4Mux_h I__10315 (
            .O(N__45502),
            .I(N__45447));
    LocalMux I__10314 (
            .O(N__45499),
            .I(N__45436));
    Span4Mux_h I__10313 (
            .O(N__45496),
            .I(N__45436));
    LocalMux I__10312 (
            .O(N__45491),
            .I(N__45436));
    LocalMux I__10311 (
            .O(N__45486),
            .I(N__45436));
    LocalMux I__10310 (
            .O(N__45483),
            .I(N__45436));
    Span4Mux_h I__10309 (
            .O(N__45478),
            .I(N__45431));
    LocalMux I__10308 (
            .O(N__45471),
            .I(N__45431));
    InMux I__10307 (
            .O(N__45470),
            .I(N__45428));
    InMux I__10306 (
            .O(N__45467),
            .I(N__45425));
    InMux I__10305 (
            .O(N__45466),
            .I(N__45420));
    InMux I__10304 (
            .O(N__45465),
            .I(N__45420));
    InMux I__10303 (
            .O(N__45464),
            .I(N__45409));
    InMux I__10302 (
            .O(N__45463),
            .I(N__45409));
    InMux I__10301 (
            .O(N__45462),
            .I(N__45409));
    InMux I__10300 (
            .O(N__45461),
            .I(N__45409));
    InMux I__10299 (
            .O(N__45460),
            .I(N__45409));
    InMux I__10298 (
            .O(N__45459),
            .I(N__45398));
    InMux I__10297 (
            .O(N__45458),
            .I(N__45398));
    InMux I__10296 (
            .O(N__45457),
            .I(N__45398));
    InMux I__10295 (
            .O(N__45456),
            .I(N__45398));
    InMux I__10294 (
            .O(N__45455),
            .I(N__45398));
    Odrv12 I__10293 (
            .O(N__45450),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk ));
    Odrv4 I__10292 (
            .O(N__45447),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk ));
    Odrv4 I__10291 (
            .O(N__45436),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk ));
    Odrv4 I__10290 (
            .O(N__45431),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk ));
    LocalMux I__10289 (
            .O(N__45428),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk ));
    LocalMux I__10288 (
            .O(N__45425),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk ));
    LocalMux I__10287 (
            .O(N__45420),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk ));
    LocalMux I__10286 (
            .O(N__45409),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk ));
    LocalMux I__10285 (
            .O(N__45398),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk ));
    CascadeMux I__10284 (
            .O(N__45379),
            .I(N__45376));
    InMux I__10283 (
            .O(N__45376),
            .I(N__45371));
    InMux I__10282 (
            .O(N__45375),
            .I(N__45365));
    InMux I__10281 (
            .O(N__45374),
            .I(N__45365));
    LocalMux I__10280 (
            .O(N__45371),
            .I(N__45361));
    InMux I__10279 (
            .O(N__45370),
            .I(N__45358));
    LocalMux I__10278 (
            .O(N__45365),
            .I(N__45355));
    CascadeMux I__10277 (
            .O(N__45364),
            .I(N__45349));
    Span4Mux_h I__10276 (
            .O(N__45361),
            .I(N__45343));
    LocalMux I__10275 (
            .O(N__45358),
            .I(N__45343));
    Span4Mux_h I__10274 (
            .O(N__45355),
            .I(N__45340));
    InMux I__10273 (
            .O(N__45354),
            .I(N__45337));
    CascadeMux I__10272 (
            .O(N__45353),
            .I(N__45329));
    CascadeMux I__10271 (
            .O(N__45352),
            .I(N__45326));
    InMux I__10270 (
            .O(N__45349),
            .I(N__45323));
    InMux I__10269 (
            .O(N__45348),
            .I(N__45320));
    Span4Mux_v I__10268 (
            .O(N__45343),
            .I(N__45317));
    Span4Mux_v I__10267 (
            .O(N__45340),
            .I(N__45306));
    LocalMux I__10266 (
            .O(N__45337),
            .I(N__45306));
    CascadeMux I__10265 (
            .O(N__45336),
            .I(N__45303));
    CascadeMux I__10264 (
            .O(N__45335),
            .I(N__45300));
    CascadeMux I__10263 (
            .O(N__45334),
            .I(N__45297));
    InMux I__10262 (
            .O(N__45333),
            .I(N__45294));
    CascadeMux I__10261 (
            .O(N__45332),
            .I(N__45291));
    InMux I__10260 (
            .O(N__45329),
            .I(N__45287));
    InMux I__10259 (
            .O(N__45326),
            .I(N__45284));
    LocalMux I__10258 (
            .O(N__45323),
            .I(N__45281));
    LocalMux I__10257 (
            .O(N__45320),
            .I(N__45276));
    Span4Mux_h I__10256 (
            .O(N__45317),
            .I(N__45276));
    InMux I__10255 (
            .O(N__45316),
            .I(N__45271));
    InMux I__10254 (
            .O(N__45315),
            .I(N__45271));
    InMux I__10253 (
            .O(N__45314),
            .I(N__45268));
    InMux I__10252 (
            .O(N__45313),
            .I(N__45265));
    InMux I__10251 (
            .O(N__45312),
            .I(N__45260));
    InMux I__10250 (
            .O(N__45311),
            .I(N__45260));
    Span4Mux_v I__10249 (
            .O(N__45306),
            .I(N__45257));
    InMux I__10248 (
            .O(N__45303),
            .I(N__45252));
    InMux I__10247 (
            .O(N__45300),
            .I(N__45252));
    InMux I__10246 (
            .O(N__45297),
            .I(N__45249));
    LocalMux I__10245 (
            .O(N__45294),
            .I(N__45246));
    InMux I__10244 (
            .O(N__45291),
            .I(N__45243));
    InMux I__10243 (
            .O(N__45290),
            .I(N__45240));
    LocalMux I__10242 (
            .O(N__45287),
            .I(N__45223));
    LocalMux I__10241 (
            .O(N__45284),
            .I(N__45223));
    Span12Mux_s11_v I__10240 (
            .O(N__45281),
            .I(N__45223));
    Sp12to4 I__10239 (
            .O(N__45276),
            .I(N__45223));
    LocalMux I__10238 (
            .O(N__45271),
            .I(N__45223));
    LocalMux I__10237 (
            .O(N__45268),
            .I(N__45223));
    LocalMux I__10236 (
            .O(N__45265),
            .I(N__45223));
    LocalMux I__10235 (
            .O(N__45260),
            .I(N__45223));
    Odrv4 I__10234 (
            .O(N__45257),
            .I(\delay_measurement_inst.delay_tr9 ));
    LocalMux I__10233 (
            .O(N__45252),
            .I(\delay_measurement_inst.delay_tr9 ));
    LocalMux I__10232 (
            .O(N__45249),
            .I(\delay_measurement_inst.delay_tr9 ));
    Odrv4 I__10231 (
            .O(N__45246),
            .I(\delay_measurement_inst.delay_tr9 ));
    LocalMux I__10230 (
            .O(N__45243),
            .I(\delay_measurement_inst.delay_tr9 ));
    LocalMux I__10229 (
            .O(N__45240),
            .I(\delay_measurement_inst.delay_tr9 ));
    Odrv12 I__10228 (
            .O(N__45223),
            .I(\delay_measurement_inst.delay_tr9 ));
    InMux I__10227 (
            .O(N__45208),
            .I(N__45205));
    LocalMux I__10226 (
            .O(N__45205),
            .I(N__45202));
    Span12Mux_v I__10225 (
            .O(N__45202),
            .I(N__45199));
    Odrv12 I__10224 (
            .O(N__45199),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ));
    InMux I__10223 (
            .O(N__45196),
            .I(N__45193));
    LocalMux I__10222 (
            .O(N__45193),
            .I(N__45190));
    Odrv4 I__10221 (
            .O(N__45190),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ));
    CascadeMux I__10220 (
            .O(N__45187),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__10219 (
            .O(N__45184),
            .I(N__45181));
    LocalMux I__10218 (
            .O(N__45181),
            .I(N__45177));
    InMux I__10217 (
            .O(N__45180),
            .I(N__45174));
    Odrv4 I__10216 (
            .O(N__45177),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__10215 (
            .O(N__45174),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    InMux I__10214 (
            .O(N__45169),
            .I(N__45165));
    InMux I__10213 (
            .O(N__45168),
            .I(N__45162));
    LocalMux I__10212 (
            .O(N__45165),
            .I(N__45159));
    LocalMux I__10211 (
            .O(N__45162),
            .I(N__45156));
    Span4Mux_h I__10210 (
            .O(N__45159),
            .I(N__45151));
    Span4Mux_h I__10209 (
            .O(N__45156),
            .I(N__45151));
    Odrv4 I__10208 (
            .O(N__45151),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__10207 (
            .O(N__45148),
            .I(N__45144));
    InMux I__10206 (
            .O(N__45147),
            .I(N__45141));
    LocalMux I__10205 (
            .O(N__45144),
            .I(N__45138));
    LocalMux I__10204 (
            .O(N__45141),
            .I(N__45135));
    Span4Mux_v I__10203 (
            .O(N__45138),
            .I(N__45130));
    Span4Mux_v I__10202 (
            .O(N__45135),
            .I(N__45130));
    Odrv4 I__10201 (
            .O(N__45130),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    CascadeMux I__10200 (
            .O(N__45127),
            .I(N__45124));
    InMux I__10199 (
            .O(N__45124),
            .I(N__45120));
    InMux I__10198 (
            .O(N__45123),
            .I(N__45117));
    LocalMux I__10197 (
            .O(N__45120),
            .I(N__45114));
    LocalMux I__10196 (
            .O(N__45117),
            .I(N__45111));
    Span4Mux_v I__10195 (
            .O(N__45114),
            .I(N__45108));
    Span4Mux_v I__10194 (
            .O(N__45111),
            .I(N__45105));
    Sp12to4 I__10193 (
            .O(N__45108),
            .I(N__45102));
    Odrv4 I__10192 (
            .O(N__45105),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv12 I__10191 (
            .O(N__45102),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__10190 (
            .O(N__45097),
            .I(N__45093));
    InMux I__10189 (
            .O(N__45096),
            .I(N__45090));
    LocalMux I__10188 (
            .O(N__45093),
            .I(N__45087));
    LocalMux I__10187 (
            .O(N__45090),
            .I(N__45084));
    Span4Mux_h I__10186 (
            .O(N__45087),
            .I(N__45081));
    Odrv4 I__10185 (
            .O(N__45084),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__10184 (
            .O(N__45081),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__10183 (
            .O(N__45076),
            .I(N__45073));
    LocalMux I__10182 (
            .O(N__45073),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19 ));
    InMux I__10181 (
            .O(N__45070),
            .I(N__45067));
    LocalMux I__10180 (
            .O(N__45067),
            .I(N__45064));
    Span4Mux_h I__10179 (
            .O(N__45064),
            .I(N__45061));
    Odrv4 I__10178 (
            .O(N__45061),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17 ));
    CascadeMux I__10177 (
            .O(N__45058),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18_cascade_ ));
    InMux I__10176 (
            .O(N__45055),
            .I(N__45052));
    LocalMux I__10175 (
            .O(N__45052),
            .I(N__45049));
    Span4Mux_v I__10174 (
            .O(N__45049),
            .I(N__45046));
    Odrv4 I__10173 (
            .O(N__45046),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16 ));
    InMux I__10172 (
            .O(N__45043),
            .I(N__45040));
    LocalMux I__10171 (
            .O(N__45040),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25 ));
    InMux I__10170 (
            .O(N__45037),
            .I(N__45034));
    LocalMux I__10169 (
            .O(N__45034),
            .I(N__45031));
    Span4Mux_h I__10168 (
            .O(N__45031),
            .I(N__45028));
    Odrv4 I__10167 (
            .O(N__45028),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df28 ));
    InMux I__10166 (
            .O(N__45025),
            .I(N__45022));
    LocalMux I__10165 (
            .O(N__45022),
            .I(N__45019));
    Span4Mux_h I__10164 (
            .O(N__45019),
            .I(N__45016));
    Odrv4 I__10163 (
            .O(N__45016),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df26 ));
    InMux I__10162 (
            .O(N__45013),
            .I(N__45010));
    LocalMux I__10161 (
            .O(N__45010),
            .I(N__45007));
    Span4Mux_v I__10160 (
            .O(N__45007),
            .I(N__45003));
    InMux I__10159 (
            .O(N__45006),
            .I(N__45000));
    Odrv4 I__10158 (
            .O(N__45003),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__10157 (
            .O(N__45000),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    CascadeMux I__10156 (
            .O(N__44995),
            .I(N__44991));
    InMux I__10155 (
            .O(N__44994),
            .I(N__44988));
    InMux I__10154 (
            .O(N__44991),
            .I(N__44984));
    LocalMux I__10153 (
            .O(N__44988),
            .I(N__44981));
    CascadeMux I__10152 (
            .O(N__44987),
            .I(N__44978));
    LocalMux I__10151 (
            .O(N__44984),
            .I(N__44975));
    Span4Mux_v I__10150 (
            .O(N__44981),
            .I(N__44972));
    InMux I__10149 (
            .O(N__44978),
            .I(N__44968));
    Span4Mux_v I__10148 (
            .O(N__44975),
            .I(N__44963));
    Span4Mux_h I__10147 (
            .O(N__44972),
            .I(N__44963));
    InMux I__10146 (
            .O(N__44971),
            .I(N__44960));
    LocalMux I__10145 (
            .O(N__44968),
            .I(elapsed_time_ns_1_RNI5GT8E1_0_13));
    Odrv4 I__10144 (
            .O(N__44963),
            .I(elapsed_time_ns_1_RNI5GT8E1_0_13));
    LocalMux I__10143 (
            .O(N__44960),
            .I(elapsed_time_ns_1_RNI5GT8E1_0_13));
    InMux I__10142 (
            .O(N__44953),
            .I(N__44950));
    LocalMux I__10141 (
            .O(N__44950),
            .I(N__44947));
    Span4Mux_h I__10140 (
            .O(N__44947),
            .I(N__44944));
    Odrv4 I__10139 (
            .O(N__44944),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ));
    CascadeMux I__10138 (
            .O(N__44941),
            .I(N__44937));
    CascadeMux I__10137 (
            .O(N__44940),
            .I(N__44934));
    InMux I__10136 (
            .O(N__44937),
            .I(N__44930));
    InMux I__10135 (
            .O(N__44934),
            .I(N__44927));
    InMux I__10134 (
            .O(N__44933),
            .I(N__44924));
    LocalMux I__10133 (
            .O(N__44930),
            .I(N__44919));
    LocalMux I__10132 (
            .O(N__44927),
            .I(N__44919));
    LocalMux I__10131 (
            .O(N__44924),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv12 I__10130 (
            .O(N__44919),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__10129 (
            .O(N__44914),
            .I(N__44911));
    LocalMux I__10128 (
            .O(N__44911),
            .I(N__44908));
    Span4Mux_h I__10127 (
            .O(N__44908),
            .I(N__44904));
    InMux I__10126 (
            .O(N__44907),
            .I(N__44901));
    Span4Mux_v I__10125 (
            .O(N__44904),
            .I(N__44898));
    LocalMux I__10124 (
            .O(N__44901),
            .I(N__44895));
    Odrv4 I__10123 (
            .O(N__44898),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__10122 (
            .O(N__44895),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__10121 (
            .O(N__44890),
            .I(bfn_17_14_0_));
    CascadeMux I__10120 (
            .O(N__44887),
            .I(N__44884));
    InMux I__10119 (
            .O(N__44884),
            .I(N__44880));
    CascadeMux I__10118 (
            .O(N__44883),
            .I(N__44877));
    LocalMux I__10117 (
            .O(N__44880),
            .I(N__44873));
    InMux I__10116 (
            .O(N__44877),
            .I(N__44870));
    InMux I__10115 (
            .O(N__44876),
            .I(N__44867));
    Sp12to4 I__10114 (
            .O(N__44873),
            .I(N__44862));
    LocalMux I__10113 (
            .O(N__44870),
            .I(N__44862));
    LocalMux I__10112 (
            .O(N__44867),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv12 I__10111 (
            .O(N__44862),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    CascadeMux I__10110 (
            .O(N__44857),
            .I(N__44854));
    InMux I__10109 (
            .O(N__44854),
            .I(N__44850));
    CascadeMux I__10108 (
            .O(N__44853),
            .I(N__44847));
    LocalMux I__10107 (
            .O(N__44850),
            .I(N__44844));
    InMux I__10106 (
            .O(N__44847),
            .I(N__44841));
    Span4Mux_h I__10105 (
            .O(N__44844),
            .I(N__44838));
    LocalMux I__10104 (
            .O(N__44841),
            .I(N__44835));
    Span4Mux_v I__10103 (
            .O(N__44838),
            .I(N__44830));
    Span4Mux_h I__10102 (
            .O(N__44835),
            .I(N__44830));
    Odrv4 I__10101 (
            .O(N__44830),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__10100 (
            .O(N__44827),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__10099 (
            .O(N__44824),
            .I(N__44820));
    InMux I__10098 (
            .O(N__44823),
            .I(N__44817));
    LocalMux I__10097 (
            .O(N__44820),
            .I(N__44814));
    LocalMux I__10096 (
            .O(N__44817),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv12 I__10095 (
            .O(N__44814),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__10094 (
            .O(N__44809),
            .I(N__44806));
    InMux I__10093 (
            .O(N__44806),
            .I(N__44801));
    InMux I__10092 (
            .O(N__44805),
            .I(N__44798));
    InMux I__10091 (
            .O(N__44804),
            .I(N__44795));
    LocalMux I__10090 (
            .O(N__44801),
            .I(N__44790));
    LocalMux I__10089 (
            .O(N__44798),
            .I(N__44790));
    LocalMux I__10088 (
            .O(N__44795),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    Odrv12 I__10087 (
            .O(N__44790),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__10086 (
            .O(N__44785),
            .I(N__44781));
    InMux I__10085 (
            .O(N__44784),
            .I(N__44778));
    LocalMux I__10084 (
            .O(N__44781),
            .I(N__44775));
    LocalMux I__10083 (
            .O(N__44778),
            .I(N__44772));
    Span4Mux_v I__10082 (
            .O(N__44775),
            .I(N__44769));
    Span4Mux_h I__10081 (
            .O(N__44772),
            .I(N__44766));
    Odrv4 I__10080 (
            .O(N__44769),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__10079 (
            .O(N__44766),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__10078 (
            .O(N__44761),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__10077 (
            .O(N__44758),
            .I(N__44753));
    InMux I__10076 (
            .O(N__44757),
            .I(N__44748));
    InMux I__10075 (
            .O(N__44756),
            .I(N__44748));
    LocalMux I__10074 (
            .O(N__44753),
            .I(N__44743));
    LocalMux I__10073 (
            .O(N__44748),
            .I(N__44743));
    Odrv12 I__10072 (
            .O(N__44743),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    CascadeMux I__10071 (
            .O(N__44740),
            .I(N__44737));
    InMux I__10070 (
            .O(N__44737),
            .I(N__44733));
    InMux I__10069 (
            .O(N__44736),
            .I(N__44730));
    LocalMux I__10068 (
            .O(N__44733),
            .I(N__44727));
    LocalMux I__10067 (
            .O(N__44730),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv12 I__10066 (
            .O(N__44727),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    InMux I__10065 (
            .O(N__44722),
            .I(N__44718));
    InMux I__10064 (
            .O(N__44721),
            .I(N__44715));
    LocalMux I__10063 (
            .O(N__44718),
            .I(N__44712));
    LocalMux I__10062 (
            .O(N__44715),
            .I(N__44709));
    Span4Mux_v I__10061 (
            .O(N__44712),
            .I(N__44704));
    Span4Mux_h I__10060 (
            .O(N__44709),
            .I(N__44704));
    Odrv4 I__10059 (
            .O(N__44704),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__10058 (
            .O(N__44701),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__10057 (
            .O(N__44698),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__10056 (
            .O(N__44695),
            .I(N__44687));
    InMux I__10055 (
            .O(N__44694),
            .I(N__44687));
    InMux I__10054 (
            .O(N__44693),
            .I(N__44684));
    CascadeMux I__10053 (
            .O(N__44692),
            .I(N__44681));
    LocalMux I__10052 (
            .O(N__44687),
            .I(N__44677));
    LocalMux I__10051 (
            .O(N__44684),
            .I(N__44674));
    InMux I__10050 (
            .O(N__44681),
            .I(N__44671));
    InMux I__10049 (
            .O(N__44680),
            .I(N__44668));
    Span4Mux_h I__10048 (
            .O(N__44677),
            .I(N__44665));
    Span4Mux_h I__10047 (
            .O(N__44674),
            .I(N__44657));
    LocalMux I__10046 (
            .O(N__44671),
            .I(N__44657));
    LocalMux I__10045 (
            .O(N__44668),
            .I(N__44657));
    Span4Mux_v I__10044 (
            .O(N__44665),
            .I(N__44654));
    InMux I__10043 (
            .O(N__44664),
            .I(N__44651));
    Span4Mux_v I__10042 (
            .O(N__44657),
            .I(N__44648));
    Odrv4 I__10041 (
            .O(N__44654),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    LocalMux I__10040 (
            .O(N__44651),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    Odrv4 I__10039 (
            .O(N__44648),
            .I(\delay_measurement_inst.elapsed_time_tr_31 ));
    InMux I__10038 (
            .O(N__44641),
            .I(N__44637));
    CascadeMux I__10037 (
            .O(N__44640),
            .I(N__44634));
    LocalMux I__10036 (
            .O(N__44637),
            .I(N__44631));
    InMux I__10035 (
            .O(N__44634),
            .I(N__44628));
    Span4Mux_h I__10034 (
            .O(N__44631),
            .I(N__44625));
    LocalMux I__10033 (
            .O(N__44628),
            .I(N__44619));
    Span4Mux_v I__10032 (
            .O(N__44625),
            .I(N__44619));
    InMux I__10031 (
            .O(N__44624),
            .I(N__44615));
    Span4Mux_v I__10030 (
            .O(N__44619),
            .I(N__44612));
    InMux I__10029 (
            .O(N__44618),
            .I(N__44609));
    LocalMux I__10028 (
            .O(N__44615),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__10027 (
            .O(N__44612),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__10026 (
            .O(N__44609),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__10025 (
            .O(N__44602),
            .I(N__44598));
    InMux I__10024 (
            .O(N__44601),
            .I(N__44594));
    LocalMux I__10023 (
            .O(N__44598),
            .I(N__44591));
    InMux I__10022 (
            .O(N__44597),
            .I(N__44588));
    LocalMux I__10021 (
            .O(N__44594),
            .I(N__44585));
    Span4Mux_v I__10020 (
            .O(N__44591),
            .I(N__44582));
    LocalMux I__10019 (
            .O(N__44588),
            .I(N__44579));
    Span4Mux_v I__10018 (
            .O(N__44585),
            .I(N__44576));
    Span4Mux_v I__10017 (
            .O(N__44582),
            .I(N__44573));
    Span4Mux_v I__10016 (
            .O(N__44579),
            .I(N__44570));
    Span4Mux_v I__10015 (
            .O(N__44576),
            .I(N__44567));
    Span4Mux_v I__10014 (
            .O(N__44573),
            .I(N__44562));
    Span4Mux_h I__10013 (
            .O(N__44570),
            .I(N__44562));
    Odrv4 I__10012 (
            .O(N__44567),
            .I(il_min_comp1_D2));
    Odrv4 I__10011 (
            .O(N__44562),
            .I(il_min_comp1_D2));
    InMux I__10010 (
            .O(N__44557),
            .I(N__44554));
    LocalMux I__10009 (
            .O(N__44554),
            .I(N__44549));
    InMux I__10008 (
            .O(N__44553),
            .I(N__44546));
    InMux I__10007 (
            .O(N__44552),
            .I(N__44543));
    Span4Mux_v I__10006 (
            .O(N__44549),
            .I(N__44536));
    LocalMux I__10005 (
            .O(N__44546),
            .I(N__44536));
    LocalMux I__10004 (
            .O(N__44543),
            .I(N__44533));
    InMux I__10003 (
            .O(N__44542),
            .I(N__44529));
    InMux I__10002 (
            .O(N__44541),
            .I(N__44526));
    Span4Mux_h I__10001 (
            .O(N__44536),
            .I(N__44523));
    Span4Mux_h I__10000 (
            .O(N__44533),
            .I(N__44520));
    InMux I__9999 (
            .O(N__44532),
            .I(N__44517));
    LocalMux I__9998 (
            .O(N__44529),
            .I(N__44512));
    LocalMux I__9997 (
            .O(N__44526),
            .I(N__44512));
    Odrv4 I__9996 (
            .O(N__44523),
            .I(phase_controller_inst1_state_4));
    Odrv4 I__9995 (
            .O(N__44520),
            .I(phase_controller_inst1_state_4));
    LocalMux I__9994 (
            .O(N__44517),
            .I(phase_controller_inst1_state_4));
    Odrv12 I__9993 (
            .O(N__44512),
            .I(phase_controller_inst1_state_4));
    InMux I__9992 (
            .O(N__44503),
            .I(N__44500));
    LocalMux I__9991 (
            .O(N__44500),
            .I(N__44497));
    Span4Mux_h I__9990 (
            .O(N__44497),
            .I(N__44494));
    Span4Mux_v I__9989 (
            .O(N__44494),
            .I(N__44491));
    Span4Mux_h I__9988 (
            .O(N__44491),
            .I(N__44487));
    InMux I__9987 (
            .O(N__44490),
            .I(N__44484));
    Odrv4 I__9986 (
            .O(N__44487),
            .I(\phase_controller_inst1.N_55 ));
    LocalMux I__9985 (
            .O(N__44484),
            .I(\phase_controller_inst1.N_55 ));
    CascadeMux I__9984 (
            .O(N__44479),
            .I(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0_cascade_ ));
    CascadeMux I__9983 (
            .O(N__44476),
            .I(N__44472));
    CascadeMux I__9982 (
            .O(N__44475),
            .I(N__44469));
    InMux I__9981 (
            .O(N__44472),
            .I(N__44466));
    InMux I__9980 (
            .O(N__44469),
            .I(N__44463));
    LocalMux I__9979 (
            .O(N__44466),
            .I(N__44457));
    LocalMux I__9978 (
            .O(N__44463),
            .I(N__44457));
    InMux I__9977 (
            .O(N__44462),
            .I(N__44454));
    Span4Mux_v I__9976 (
            .O(N__44457),
            .I(N__44451));
    LocalMux I__9975 (
            .O(N__44454),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__9974 (
            .O(N__44451),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__9973 (
            .O(N__44446),
            .I(bfn_17_13_0_));
    CascadeMux I__9972 (
            .O(N__44443),
            .I(N__44440));
    InMux I__9971 (
            .O(N__44440),
            .I(N__44437));
    LocalMux I__9970 (
            .O(N__44437),
            .I(N__44432));
    InMux I__9969 (
            .O(N__44436),
            .I(N__44429));
    InMux I__9968 (
            .O(N__44435),
            .I(N__44426));
    Sp12to4 I__9967 (
            .O(N__44432),
            .I(N__44421));
    LocalMux I__9966 (
            .O(N__44429),
            .I(N__44421));
    LocalMux I__9965 (
            .O(N__44426),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv12 I__9964 (
            .O(N__44421),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__9963 (
            .O(N__44416),
            .I(N__44413));
    LocalMux I__9962 (
            .O(N__44413),
            .I(N__44410));
    Span4Mux_v I__9961 (
            .O(N__44410),
            .I(N__44406));
    InMux I__9960 (
            .O(N__44409),
            .I(N__44403));
    Odrv4 I__9959 (
            .O(N__44406),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__9958 (
            .O(N__44403),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__9957 (
            .O(N__44398),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__9956 (
            .O(N__44395),
            .I(N__44388));
    InMux I__9955 (
            .O(N__44394),
            .I(N__44388));
    InMux I__9954 (
            .O(N__44393),
            .I(N__44385));
    LocalMux I__9953 (
            .O(N__44388),
            .I(N__44382));
    LocalMux I__9952 (
            .O(N__44385),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    Odrv12 I__9951 (
            .O(N__44382),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__9950 (
            .O(N__44377),
            .I(N__44374));
    LocalMux I__9949 (
            .O(N__44374),
            .I(N__44371));
    Span4Mux_h I__9948 (
            .O(N__44371),
            .I(N__44367));
    InMux I__9947 (
            .O(N__44370),
            .I(N__44364));
    Odrv4 I__9946 (
            .O(N__44367),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__9945 (
            .O(N__44364),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__9944 (
            .O(N__44359),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__9943 (
            .O(N__44356),
            .I(N__44349));
    InMux I__9942 (
            .O(N__44355),
            .I(N__44349));
    InMux I__9941 (
            .O(N__44354),
            .I(N__44346));
    LocalMux I__9940 (
            .O(N__44349),
            .I(N__44343));
    LocalMux I__9939 (
            .O(N__44346),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv12 I__9938 (
            .O(N__44343),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__9937 (
            .O(N__44338),
            .I(N__44335));
    LocalMux I__9936 (
            .O(N__44335),
            .I(N__44332));
    Span4Mux_h I__9935 (
            .O(N__44332),
            .I(N__44328));
    InMux I__9934 (
            .O(N__44331),
            .I(N__44325));
    Odrv4 I__9933 (
            .O(N__44328),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    LocalMux I__9932 (
            .O(N__44325),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__9931 (
            .O(N__44320),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__9930 (
            .O(N__44317),
            .I(N__44313));
    CascadeMux I__9929 (
            .O(N__44316),
            .I(N__44310));
    InMux I__9928 (
            .O(N__44313),
            .I(N__44304));
    InMux I__9927 (
            .O(N__44310),
            .I(N__44304));
    InMux I__9926 (
            .O(N__44309),
            .I(N__44301));
    LocalMux I__9925 (
            .O(N__44304),
            .I(N__44298));
    LocalMux I__9924 (
            .O(N__44301),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv12 I__9923 (
            .O(N__44298),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__9922 (
            .O(N__44293),
            .I(N__44290));
    LocalMux I__9921 (
            .O(N__44290),
            .I(N__44286));
    InMux I__9920 (
            .O(N__44289),
            .I(N__44283));
    Span4Mux_v I__9919 (
            .O(N__44286),
            .I(N__44278));
    LocalMux I__9918 (
            .O(N__44283),
            .I(N__44278));
    Odrv4 I__9917 (
            .O(N__44278),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__9916 (
            .O(N__44275),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__9915 (
            .O(N__44272),
            .I(N__44268));
    CascadeMux I__9914 (
            .O(N__44271),
            .I(N__44265));
    InMux I__9913 (
            .O(N__44268),
            .I(N__44259));
    InMux I__9912 (
            .O(N__44265),
            .I(N__44259));
    InMux I__9911 (
            .O(N__44264),
            .I(N__44256));
    LocalMux I__9910 (
            .O(N__44259),
            .I(N__44253));
    LocalMux I__9909 (
            .O(N__44256),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv12 I__9908 (
            .O(N__44253),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__9907 (
            .O(N__44248),
            .I(N__44245));
    LocalMux I__9906 (
            .O(N__44245),
            .I(N__44241));
    InMux I__9905 (
            .O(N__44244),
            .I(N__44238));
    Span4Mux_h I__9904 (
            .O(N__44241),
            .I(N__44233));
    LocalMux I__9903 (
            .O(N__44238),
            .I(N__44233));
    Odrv4 I__9902 (
            .O(N__44233),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__9901 (
            .O(N__44230),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__9900 (
            .O(N__44227),
            .I(N__44221));
    InMux I__9899 (
            .O(N__44226),
            .I(N__44221));
    LocalMux I__9898 (
            .O(N__44221),
            .I(N__44217));
    InMux I__9897 (
            .O(N__44220),
            .I(N__44214));
    Span4Mux_v I__9896 (
            .O(N__44217),
            .I(N__44211));
    LocalMux I__9895 (
            .O(N__44214),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv4 I__9894 (
            .O(N__44211),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    CascadeMux I__9893 (
            .O(N__44206),
            .I(N__44203));
    InMux I__9892 (
            .O(N__44203),
            .I(N__44200));
    LocalMux I__9891 (
            .O(N__44200),
            .I(N__44197));
    Span12Mux_v I__9890 (
            .O(N__44197),
            .I(N__44193));
    InMux I__9889 (
            .O(N__44196),
            .I(N__44190));
    Odrv12 I__9888 (
            .O(N__44193),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__9887 (
            .O(N__44190),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__9886 (
            .O(N__44185),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__9885 (
            .O(N__44182),
            .I(N__44176));
    InMux I__9884 (
            .O(N__44181),
            .I(N__44176));
    LocalMux I__9883 (
            .O(N__44176),
            .I(N__44172));
    InMux I__9882 (
            .O(N__44175),
            .I(N__44169));
    Span4Mux_v I__9881 (
            .O(N__44172),
            .I(N__44166));
    LocalMux I__9880 (
            .O(N__44169),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__9879 (
            .O(N__44166),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__9878 (
            .O(N__44161),
            .I(N__44158));
    LocalMux I__9877 (
            .O(N__44158),
            .I(N__44154));
    InMux I__9876 (
            .O(N__44157),
            .I(N__44151));
    Span4Mux_h I__9875 (
            .O(N__44154),
            .I(N__44148));
    LocalMux I__9874 (
            .O(N__44151),
            .I(N__44145));
    Span4Mux_v I__9873 (
            .O(N__44148),
            .I(N__44142));
    Span4Mux_h I__9872 (
            .O(N__44145),
            .I(N__44139));
    Odrv4 I__9871 (
            .O(N__44142),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv4 I__9870 (
            .O(N__44139),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__9869 (
            .O(N__44134),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__9868 (
            .O(N__44131),
            .I(N__44128));
    InMux I__9867 (
            .O(N__44128),
            .I(N__44124));
    CascadeMux I__9866 (
            .O(N__44127),
            .I(N__44121));
    LocalMux I__9865 (
            .O(N__44124),
            .I(N__44117));
    InMux I__9864 (
            .O(N__44121),
            .I(N__44114));
    InMux I__9863 (
            .O(N__44120),
            .I(N__44111));
    Sp12to4 I__9862 (
            .O(N__44117),
            .I(N__44106));
    LocalMux I__9861 (
            .O(N__44114),
            .I(N__44106));
    LocalMux I__9860 (
            .O(N__44111),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv12 I__9859 (
            .O(N__44106),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__9858 (
            .O(N__44101),
            .I(N__44098));
    LocalMux I__9857 (
            .O(N__44098),
            .I(N__44095));
    Span4Mux_v I__9856 (
            .O(N__44095),
            .I(N__44091));
    InMux I__9855 (
            .O(N__44094),
            .I(N__44088));
    Odrv4 I__9854 (
            .O(N__44091),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__9853 (
            .O(N__44088),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__9852 (
            .O(N__44083),
            .I(bfn_17_12_0_));
    CascadeMux I__9851 (
            .O(N__44080),
            .I(N__44076));
    CascadeMux I__9850 (
            .O(N__44079),
            .I(N__44073));
    InMux I__9849 (
            .O(N__44076),
            .I(N__44069));
    InMux I__9848 (
            .O(N__44073),
            .I(N__44066));
    InMux I__9847 (
            .O(N__44072),
            .I(N__44063));
    LocalMux I__9846 (
            .O(N__44069),
            .I(N__44058));
    LocalMux I__9845 (
            .O(N__44066),
            .I(N__44058));
    LocalMux I__9844 (
            .O(N__44063),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    Odrv12 I__9843 (
            .O(N__44058),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__9842 (
            .O(N__44053),
            .I(N__44050));
    LocalMux I__9841 (
            .O(N__44050),
            .I(N__44047));
    Span4Mux_h I__9840 (
            .O(N__44047),
            .I(N__44043));
    InMux I__9839 (
            .O(N__44046),
            .I(N__44040));
    Odrv4 I__9838 (
            .O(N__44043),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    LocalMux I__9837 (
            .O(N__44040),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__9836 (
            .O(N__44035),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__9835 (
            .O(N__44032),
            .I(N__44026));
    InMux I__9834 (
            .O(N__44031),
            .I(N__44026));
    LocalMux I__9833 (
            .O(N__44026),
            .I(N__44022));
    InMux I__9832 (
            .O(N__44025),
            .I(N__44019));
    Span4Mux_v I__9831 (
            .O(N__44022),
            .I(N__44016));
    LocalMux I__9830 (
            .O(N__44019),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__9829 (
            .O(N__44016),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__9828 (
            .O(N__44011),
            .I(N__44008));
    LocalMux I__9827 (
            .O(N__44008),
            .I(N__44004));
    CascadeMux I__9826 (
            .O(N__44007),
            .I(N__44001));
    Span4Mux_v I__9825 (
            .O(N__44004),
            .I(N__43998));
    InMux I__9824 (
            .O(N__44001),
            .I(N__43995));
    Odrv4 I__9823 (
            .O(N__43998),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__9822 (
            .O(N__43995),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__9821 (
            .O(N__43990),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__9820 (
            .O(N__43987),
            .I(N__43984));
    InMux I__9819 (
            .O(N__43984),
            .I(N__43981));
    LocalMux I__9818 (
            .O(N__43981),
            .I(N__43977));
    InMux I__9817 (
            .O(N__43980),
            .I(N__43974));
    Span4Mux_h I__9816 (
            .O(N__43977),
            .I(N__43968));
    LocalMux I__9815 (
            .O(N__43974),
            .I(N__43968));
    InMux I__9814 (
            .O(N__43973),
            .I(N__43965));
    Span4Mux_v I__9813 (
            .O(N__43968),
            .I(N__43962));
    LocalMux I__9812 (
            .O(N__43965),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv4 I__9811 (
            .O(N__43962),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__9810 (
            .O(N__43957),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__9809 (
            .O(N__43954),
            .I(N__43950));
    CascadeMux I__9808 (
            .O(N__43953),
            .I(N__43947));
    InMux I__9807 (
            .O(N__43950),
            .I(N__43941));
    InMux I__9806 (
            .O(N__43947),
            .I(N__43941));
    InMux I__9805 (
            .O(N__43946),
            .I(N__43938));
    LocalMux I__9804 (
            .O(N__43941),
            .I(N__43935));
    LocalMux I__9803 (
            .O(N__43938),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv12 I__9802 (
            .O(N__43935),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__9801 (
            .O(N__43930),
            .I(N__43926));
    InMux I__9800 (
            .O(N__43929),
            .I(N__43923));
    LocalMux I__9799 (
            .O(N__43926),
            .I(N__43920));
    LocalMux I__9798 (
            .O(N__43923),
            .I(N__43917));
    Span4Mux_h I__9797 (
            .O(N__43920),
            .I(N__43911));
    Span4Mux_v I__9796 (
            .O(N__43917),
            .I(N__43911));
    InMux I__9795 (
            .O(N__43916),
            .I(N__43908));
    Odrv4 I__9794 (
            .O(N__43911),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    LocalMux I__9793 (
            .O(N__43908),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ));
    InMux I__9792 (
            .O(N__43903),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__9791 (
            .O(N__43900),
            .I(N__43893));
    InMux I__9790 (
            .O(N__43899),
            .I(N__43893));
    InMux I__9789 (
            .O(N__43898),
            .I(N__43890));
    LocalMux I__9788 (
            .O(N__43893),
            .I(N__43887));
    LocalMux I__9787 (
            .O(N__43890),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv12 I__9786 (
            .O(N__43887),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__9785 (
            .O(N__43882),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__9784 (
            .O(N__43879),
            .I(N__43873));
    InMux I__9783 (
            .O(N__43878),
            .I(N__43873));
    LocalMux I__9782 (
            .O(N__43873),
            .I(N__43869));
    InMux I__9781 (
            .O(N__43872),
            .I(N__43866));
    Span4Mux_v I__9780 (
            .O(N__43869),
            .I(N__43863));
    LocalMux I__9779 (
            .O(N__43866),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv4 I__9778 (
            .O(N__43863),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__9777 (
            .O(N__43858),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__9776 (
            .O(N__43855),
            .I(N__43851));
    CascadeMux I__9775 (
            .O(N__43854),
            .I(N__43848));
    InMux I__9774 (
            .O(N__43851),
            .I(N__43843));
    InMux I__9773 (
            .O(N__43848),
            .I(N__43843));
    LocalMux I__9772 (
            .O(N__43843),
            .I(N__43839));
    InMux I__9771 (
            .O(N__43842),
            .I(N__43836));
    Span4Mux_v I__9770 (
            .O(N__43839),
            .I(N__43833));
    LocalMux I__9769 (
            .O(N__43836),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    Odrv4 I__9768 (
            .O(N__43833),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__9767 (
            .O(N__43828),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__9766 (
            .O(N__43825),
            .I(N__43799));
    InMux I__9765 (
            .O(N__43824),
            .I(N__43799));
    InMux I__9764 (
            .O(N__43823),
            .I(N__43799));
    InMux I__9763 (
            .O(N__43822),
            .I(N__43799));
    InMux I__9762 (
            .O(N__43821),
            .I(N__43790));
    InMux I__9761 (
            .O(N__43820),
            .I(N__43790));
    InMux I__9760 (
            .O(N__43819),
            .I(N__43790));
    InMux I__9759 (
            .O(N__43818),
            .I(N__43790));
    InMux I__9758 (
            .O(N__43817),
            .I(N__43781));
    InMux I__9757 (
            .O(N__43816),
            .I(N__43781));
    InMux I__9756 (
            .O(N__43815),
            .I(N__43781));
    InMux I__9755 (
            .O(N__43814),
            .I(N__43781));
    InMux I__9754 (
            .O(N__43813),
            .I(N__43764));
    InMux I__9753 (
            .O(N__43812),
            .I(N__43764));
    InMux I__9752 (
            .O(N__43811),
            .I(N__43755));
    InMux I__9751 (
            .O(N__43810),
            .I(N__43755));
    InMux I__9750 (
            .O(N__43809),
            .I(N__43755));
    InMux I__9749 (
            .O(N__43808),
            .I(N__43755));
    LocalMux I__9748 (
            .O(N__43799),
            .I(N__43748));
    LocalMux I__9747 (
            .O(N__43790),
            .I(N__43748));
    LocalMux I__9746 (
            .O(N__43781),
            .I(N__43748));
    InMux I__9745 (
            .O(N__43780),
            .I(N__43739));
    InMux I__9744 (
            .O(N__43779),
            .I(N__43739));
    InMux I__9743 (
            .O(N__43778),
            .I(N__43739));
    InMux I__9742 (
            .O(N__43777),
            .I(N__43739));
    InMux I__9741 (
            .O(N__43776),
            .I(N__43730));
    InMux I__9740 (
            .O(N__43775),
            .I(N__43730));
    InMux I__9739 (
            .O(N__43774),
            .I(N__43730));
    InMux I__9738 (
            .O(N__43773),
            .I(N__43730));
    InMux I__9737 (
            .O(N__43772),
            .I(N__43721));
    InMux I__9736 (
            .O(N__43771),
            .I(N__43721));
    InMux I__9735 (
            .O(N__43770),
            .I(N__43721));
    InMux I__9734 (
            .O(N__43769),
            .I(N__43721));
    LocalMux I__9733 (
            .O(N__43764),
            .I(N__43718));
    LocalMux I__9732 (
            .O(N__43755),
            .I(N__43715));
    Span4Mux_v I__9731 (
            .O(N__43748),
            .I(N__43710));
    LocalMux I__9730 (
            .O(N__43739),
            .I(N__43710));
    LocalMux I__9729 (
            .O(N__43730),
            .I(N__43705));
    LocalMux I__9728 (
            .O(N__43721),
            .I(N__43705));
    Span4Mux_h I__9727 (
            .O(N__43718),
            .I(N__43700));
    Span4Mux_h I__9726 (
            .O(N__43715),
            .I(N__43700));
    Span4Mux_h I__9725 (
            .O(N__43710),
            .I(N__43697));
    Odrv4 I__9724 (
            .O(N__43705),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__9723 (
            .O(N__43700),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__9722 (
            .O(N__43697),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__9721 (
            .O(N__43690),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__9720 (
            .O(N__43687),
            .I(N__43684));
    LocalMux I__9719 (
            .O(N__43684),
            .I(N__43680));
    CEMux I__9718 (
            .O(N__43683),
            .I(N__43677));
    Span4Mux_h I__9717 (
            .O(N__43680),
            .I(N__43670));
    LocalMux I__9716 (
            .O(N__43677),
            .I(N__43670));
    CEMux I__9715 (
            .O(N__43676),
            .I(N__43667));
    CEMux I__9714 (
            .O(N__43675),
            .I(N__43664));
    Span4Mux_v I__9713 (
            .O(N__43670),
            .I(N__43661));
    LocalMux I__9712 (
            .O(N__43667),
            .I(N__43658));
    LocalMux I__9711 (
            .O(N__43664),
            .I(N__43655));
    Span4Mux_h I__9710 (
            .O(N__43661),
            .I(N__43652));
    Span4Mux_h I__9709 (
            .O(N__43658),
            .I(N__43649));
    Span4Mux_h I__9708 (
            .O(N__43655),
            .I(N__43646));
    Span4Mux_h I__9707 (
            .O(N__43652),
            .I(N__43643));
    Span4Mux_h I__9706 (
            .O(N__43649),
            .I(N__43640));
    Span4Mux_h I__9705 (
            .O(N__43646),
            .I(N__43637));
    Odrv4 I__9704 (
            .O(N__43643),
            .I(\delay_measurement_inst.delay_tr_timer.N_400_i ));
    Odrv4 I__9703 (
            .O(N__43640),
            .I(\delay_measurement_inst.delay_tr_timer.N_400_i ));
    Odrv4 I__9702 (
            .O(N__43637),
            .I(\delay_measurement_inst.delay_tr_timer.N_400_i ));
    InMux I__9701 (
            .O(N__43630),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__9700 (
            .O(N__43627),
            .I(N__43621));
    InMux I__9699 (
            .O(N__43626),
            .I(N__43621));
    LocalMux I__9698 (
            .O(N__43621),
            .I(N__43617));
    InMux I__9697 (
            .O(N__43620),
            .I(N__43614));
    Span4Mux_v I__9696 (
            .O(N__43617),
            .I(N__43611));
    LocalMux I__9695 (
            .O(N__43614),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv4 I__9694 (
            .O(N__43611),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__9693 (
            .O(N__43606),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__9692 (
            .O(N__43603),
            .I(N__43597));
    InMux I__9691 (
            .O(N__43602),
            .I(N__43597));
    LocalMux I__9690 (
            .O(N__43597),
            .I(N__43593));
    InMux I__9689 (
            .O(N__43596),
            .I(N__43590));
    Span4Mux_v I__9688 (
            .O(N__43593),
            .I(N__43587));
    LocalMux I__9687 (
            .O(N__43590),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__9686 (
            .O(N__43587),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__9685 (
            .O(N__43582),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__9684 (
            .O(N__43579),
            .I(N__43575));
    CascadeMux I__9683 (
            .O(N__43578),
            .I(N__43572));
    InMux I__9682 (
            .O(N__43575),
            .I(N__43566));
    InMux I__9681 (
            .O(N__43572),
            .I(N__43566));
    InMux I__9680 (
            .O(N__43571),
            .I(N__43563));
    LocalMux I__9679 (
            .O(N__43566),
            .I(N__43560));
    LocalMux I__9678 (
            .O(N__43563),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv12 I__9677 (
            .O(N__43560),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__9676 (
            .O(N__43555),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__9675 (
            .O(N__43552),
            .I(N__43548));
    CascadeMux I__9674 (
            .O(N__43551),
            .I(N__43545));
    InMux I__9673 (
            .O(N__43548),
            .I(N__43539));
    InMux I__9672 (
            .O(N__43545),
            .I(N__43539));
    InMux I__9671 (
            .O(N__43544),
            .I(N__43536));
    LocalMux I__9670 (
            .O(N__43539),
            .I(N__43533));
    LocalMux I__9669 (
            .O(N__43536),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv12 I__9668 (
            .O(N__43533),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__9667 (
            .O(N__43528),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__9666 (
            .O(N__43525),
            .I(N__43519));
    InMux I__9665 (
            .O(N__43524),
            .I(N__43519));
    LocalMux I__9664 (
            .O(N__43519),
            .I(N__43515));
    InMux I__9663 (
            .O(N__43518),
            .I(N__43512));
    Span4Mux_v I__9662 (
            .O(N__43515),
            .I(N__43509));
    LocalMux I__9661 (
            .O(N__43512),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    Odrv4 I__9660 (
            .O(N__43509),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__9659 (
            .O(N__43504),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__9658 (
            .O(N__43501),
            .I(N__43495));
    InMux I__9657 (
            .O(N__43500),
            .I(N__43495));
    LocalMux I__9656 (
            .O(N__43495),
            .I(N__43491));
    InMux I__9655 (
            .O(N__43494),
            .I(N__43488));
    Span4Mux_v I__9654 (
            .O(N__43491),
            .I(N__43485));
    LocalMux I__9653 (
            .O(N__43488),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv4 I__9652 (
            .O(N__43485),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__9651 (
            .O(N__43480),
            .I(N__43477));
    LocalMux I__9650 (
            .O(N__43477),
            .I(N__43473));
    InMux I__9649 (
            .O(N__43476),
            .I(N__43470));
    Odrv12 I__9648 (
            .O(N__43473),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__9647 (
            .O(N__43470),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__9646 (
            .O(N__43465),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__9645 (
            .O(N__43462),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__9644 (
            .O(N__43459),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__9643 (
            .O(N__43456),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__9642 (
            .O(N__43453),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__9641 (
            .O(N__43450),
            .I(bfn_17_10_0_));
    InMux I__9640 (
            .O(N__43447),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__9639 (
            .O(N__43444),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__9638 (
            .O(N__43441),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__9637 (
            .O(N__43438),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__9636 (
            .O(N__43435),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__9635 (
            .O(N__43432),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__9634 (
            .O(N__43429),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__9633 (
            .O(N__43426),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__9632 (
            .O(N__43423),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__9631 (
            .O(N__43420),
            .I(bfn_17_9_0_));
    InMux I__9630 (
            .O(N__43417),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__9629 (
            .O(N__43414),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__9628 (
            .O(N__43411),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__9627 (
            .O(N__43408),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__9626 (
            .O(N__43405),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__9625 (
            .O(N__43402),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__9624 (
            .O(N__43399),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__9623 (
            .O(N__43396),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__9622 (
            .O(N__43393),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__9621 (
            .O(N__43390),
            .I(bfn_17_8_0_));
    InMux I__9620 (
            .O(N__43387),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__9619 (
            .O(N__43384),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    CascadeMux I__9618 (
            .O(N__43381),
            .I(N__43378));
    InMux I__9617 (
            .O(N__43378),
            .I(N__43372));
    InMux I__9616 (
            .O(N__43377),
            .I(N__43369));
    CascadeMux I__9615 (
            .O(N__43376),
            .I(N__43366));
    InMux I__9614 (
            .O(N__43375),
            .I(N__43363));
    LocalMux I__9613 (
            .O(N__43372),
            .I(N__43358));
    LocalMux I__9612 (
            .O(N__43369),
            .I(N__43358));
    InMux I__9611 (
            .O(N__43366),
            .I(N__43355));
    LocalMux I__9610 (
            .O(N__43363),
            .I(N__43352));
    Odrv12 I__9609 (
            .O(N__43358),
            .I(elapsed_time_ns_1_RNIHHC6P1_0_18));
    LocalMux I__9608 (
            .O(N__43355),
            .I(elapsed_time_ns_1_RNIHHC6P1_0_18));
    Odrv4 I__9607 (
            .O(N__43352),
            .I(elapsed_time_ns_1_RNIHHC6P1_0_18));
    InMux I__9606 (
            .O(N__43345),
            .I(N__43341));
    CascadeMux I__9605 (
            .O(N__43344),
            .I(N__43338));
    LocalMux I__9604 (
            .O(N__43341),
            .I(N__43335));
    InMux I__9603 (
            .O(N__43338),
            .I(N__43332));
    Span12Mux_s8_v I__9602 (
            .O(N__43335),
            .I(N__43329));
    LocalMux I__9601 (
            .O(N__43332),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    Odrv12 I__9600 (
            .O(N__43329),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    InMux I__9599 (
            .O(N__43324),
            .I(N__43321));
    LocalMux I__9598 (
            .O(N__43321),
            .I(N__43318));
    Span4Mux_h I__9597 (
            .O(N__43318),
            .I(N__43315));
    Span4Mux_h I__9596 (
            .O(N__43315),
            .I(N__43312));
    Odrv4 I__9595 (
            .O(N__43312),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__9594 (
            .O(N__43309),
            .I(N__43305));
    InMux I__9593 (
            .O(N__43308),
            .I(N__43302));
    InMux I__9592 (
            .O(N__43305),
            .I(N__43299));
    LocalMux I__9591 (
            .O(N__43302),
            .I(N__43292));
    LocalMux I__9590 (
            .O(N__43299),
            .I(N__43292));
    InMux I__9589 (
            .O(N__43298),
            .I(N__43289));
    InMux I__9588 (
            .O(N__43297),
            .I(N__43286));
    Span4Mux_v I__9587 (
            .O(N__43292),
            .I(N__43281));
    LocalMux I__9586 (
            .O(N__43289),
            .I(N__43281));
    LocalMux I__9585 (
            .O(N__43286),
            .I(elapsed_time_ns_1_RNI2DT8E1_0_10));
    Odrv4 I__9584 (
            .O(N__43281),
            .I(elapsed_time_ns_1_RNI2DT8E1_0_10));
    InMux I__9583 (
            .O(N__43276),
            .I(N__43273));
    LocalMux I__9582 (
            .O(N__43273),
            .I(N__43270));
    Span12Mux_h I__9581 (
            .O(N__43270),
            .I(N__43267));
    Odrv12 I__9580 (
            .O(N__43267),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__9579 (
            .O(N__43264),
            .I(N__43260));
    InMux I__9578 (
            .O(N__43263),
            .I(N__43256));
    InMux I__9577 (
            .O(N__43260),
            .I(N__43253));
    CascadeMux I__9576 (
            .O(N__43259),
            .I(N__43250));
    LocalMux I__9575 (
            .O(N__43256),
            .I(N__43244));
    LocalMux I__9574 (
            .O(N__43253),
            .I(N__43244));
    InMux I__9573 (
            .O(N__43250),
            .I(N__43239));
    InMux I__9572 (
            .O(N__43249),
            .I(N__43239));
    Odrv12 I__9571 (
            .O(N__43244),
            .I(elapsed_time_ns_1_RNI3ET8E1_0_11));
    LocalMux I__9570 (
            .O(N__43239),
            .I(elapsed_time_ns_1_RNI3ET8E1_0_11));
    InMux I__9569 (
            .O(N__43234),
            .I(N__43231));
    LocalMux I__9568 (
            .O(N__43231),
            .I(N__43228));
    Span4Mux_h I__9567 (
            .O(N__43228),
            .I(N__43225));
    Span4Mux_h I__9566 (
            .O(N__43225),
            .I(N__43222));
    Odrv4 I__9565 (
            .O(N__43222),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    CascadeMux I__9564 (
            .O(N__43219),
            .I(N__43216));
    InMux I__9563 (
            .O(N__43216),
            .I(N__43212));
    InMux I__9562 (
            .O(N__43215),
            .I(N__43209));
    LocalMux I__9561 (
            .O(N__43212),
            .I(N__43203));
    LocalMux I__9560 (
            .O(N__43209),
            .I(N__43203));
    InMux I__9559 (
            .O(N__43208),
            .I(N__43200));
    Odrv12 I__9558 (
            .O(N__43203),
            .I(elapsed_time_ns_1_RNI4FT8E1_0_12));
    LocalMux I__9557 (
            .O(N__43200),
            .I(elapsed_time_ns_1_RNI4FT8E1_0_12));
    InMux I__9556 (
            .O(N__43195),
            .I(N__43192));
    LocalMux I__9555 (
            .O(N__43192),
            .I(N__43189));
    Span4Mux_h I__9554 (
            .O(N__43189),
            .I(N__43186));
    Span4Mux_h I__9553 (
            .O(N__43186),
            .I(N__43183));
    Odrv4 I__9552 (
            .O(N__43183),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__9551 (
            .O(N__43180),
            .I(N__43177));
    LocalMux I__9550 (
            .O(N__43177),
            .I(N__43174));
    Span4Mux_h I__9549 (
            .O(N__43174),
            .I(N__43171));
    Span4Mux_h I__9548 (
            .O(N__43171),
            .I(N__43168));
    Odrv4 I__9547 (
            .O(N__43168),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__9546 (
            .O(N__43165),
            .I(N__43162));
    LocalMux I__9545 (
            .O(N__43162),
            .I(N__43159));
    Span4Mux_h I__9544 (
            .O(N__43159),
            .I(N__43156));
    Span4Mux_h I__9543 (
            .O(N__43156),
            .I(N__43153));
    Odrv4 I__9542 (
            .O(N__43153),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    CEMux I__9541 (
            .O(N__43150),
            .I(N__43145));
    CEMux I__9540 (
            .O(N__43149),
            .I(N__43118));
    CEMux I__9539 (
            .O(N__43148),
            .I(N__43115));
    LocalMux I__9538 (
            .O(N__43145),
            .I(N__43112));
    CEMux I__9537 (
            .O(N__43144),
            .I(N__43109));
    CEMux I__9536 (
            .O(N__43143),
            .I(N__43106));
    InMux I__9535 (
            .O(N__43142),
            .I(N__43097));
    InMux I__9534 (
            .O(N__43141),
            .I(N__43097));
    InMux I__9533 (
            .O(N__43140),
            .I(N__43097));
    InMux I__9532 (
            .O(N__43139),
            .I(N__43097));
    InMux I__9531 (
            .O(N__43138),
            .I(N__43082));
    InMux I__9530 (
            .O(N__43137),
            .I(N__43082));
    InMux I__9529 (
            .O(N__43136),
            .I(N__43082));
    InMux I__9528 (
            .O(N__43135),
            .I(N__43073));
    InMux I__9527 (
            .O(N__43134),
            .I(N__43073));
    InMux I__9526 (
            .O(N__43133),
            .I(N__43073));
    InMux I__9525 (
            .O(N__43132),
            .I(N__43073));
    InMux I__9524 (
            .O(N__43131),
            .I(N__43064));
    InMux I__9523 (
            .O(N__43130),
            .I(N__43064));
    InMux I__9522 (
            .O(N__43129),
            .I(N__43064));
    InMux I__9521 (
            .O(N__43128),
            .I(N__43064));
    InMux I__9520 (
            .O(N__43127),
            .I(N__43055));
    InMux I__9519 (
            .O(N__43126),
            .I(N__43055));
    InMux I__9518 (
            .O(N__43125),
            .I(N__43055));
    InMux I__9517 (
            .O(N__43124),
            .I(N__43055));
    InMux I__9516 (
            .O(N__43123),
            .I(N__43048));
    InMux I__9515 (
            .O(N__43122),
            .I(N__43048));
    InMux I__9514 (
            .O(N__43121),
            .I(N__43048));
    LocalMux I__9513 (
            .O(N__43118),
            .I(N__43043));
    LocalMux I__9512 (
            .O(N__43115),
            .I(N__43043));
    Span4Mux_v I__9511 (
            .O(N__43112),
            .I(N__43037));
    LocalMux I__9510 (
            .O(N__43109),
            .I(N__43037));
    LocalMux I__9509 (
            .O(N__43106),
            .I(N__43034));
    LocalMux I__9508 (
            .O(N__43097),
            .I(N__43031));
    InMux I__9507 (
            .O(N__43096),
            .I(N__43022));
    InMux I__9506 (
            .O(N__43095),
            .I(N__43022));
    InMux I__9505 (
            .O(N__43094),
            .I(N__43022));
    InMux I__9504 (
            .O(N__43093),
            .I(N__43022));
    InMux I__9503 (
            .O(N__43092),
            .I(N__43013));
    InMux I__9502 (
            .O(N__43091),
            .I(N__43013));
    InMux I__9501 (
            .O(N__43090),
            .I(N__43013));
    InMux I__9500 (
            .O(N__43089),
            .I(N__43013));
    LocalMux I__9499 (
            .O(N__43082),
            .I(N__43006));
    LocalMux I__9498 (
            .O(N__43073),
            .I(N__43006));
    LocalMux I__9497 (
            .O(N__43064),
            .I(N__43006));
    LocalMux I__9496 (
            .O(N__43055),
            .I(N__43001));
    LocalMux I__9495 (
            .O(N__43048),
            .I(N__43001));
    Span4Mux_v I__9494 (
            .O(N__43043),
            .I(N__42998));
    InMux I__9493 (
            .O(N__43042),
            .I(N__42995));
    Span4Mux_h I__9492 (
            .O(N__43037),
            .I(N__42992));
    Span4Mux_v I__9491 (
            .O(N__43034),
            .I(N__42979));
    Span4Mux_v I__9490 (
            .O(N__43031),
            .I(N__42979));
    LocalMux I__9489 (
            .O(N__43022),
            .I(N__42979));
    LocalMux I__9488 (
            .O(N__43013),
            .I(N__42979));
    Span4Mux_v I__9487 (
            .O(N__43006),
            .I(N__42979));
    Span4Mux_v I__9486 (
            .O(N__43001),
            .I(N__42979));
    Odrv4 I__9485 (
            .O(N__42998),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__9484 (
            .O(N__42995),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__9483 (
            .O(N__42992),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__9482 (
            .O(N__42979),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__9481 (
            .O(N__42970),
            .I(bfn_17_7_0_));
    InMux I__9480 (
            .O(N__42967),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__9479 (
            .O(N__42964),
            .I(N__42959));
    InMux I__9478 (
            .O(N__42963),
            .I(N__42956));
    InMux I__9477 (
            .O(N__42962),
            .I(N__42951));
    LocalMux I__9476 (
            .O(N__42959),
            .I(N__42946));
    LocalMux I__9475 (
            .O(N__42956),
            .I(N__42946));
    InMux I__9474 (
            .O(N__42955),
            .I(N__42943));
    InMux I__9473 (
            .O(N__42954),
            .I(N__42940));
    LocalMux I__9472 (
            .O(N__42951),
            .I(elapsed_time_ns_1_RNIIIC6P1_0_19));
    Odrv12 I__9471 (
            .O(N__42946),
            .I(elapsed_time_ns_1_RNIIIC6P1_0_19));
    LocalMux I__9470 (
            .O(N__42943),
            .I(elapsed_time_ns_1_RNIIIC6P1_0_19));
    LocalMux I__9469 (
            .O(N__42940),
            .I(elapsed_time_ns_1_RNIIIC6P1_0_19));
    CascadeMux I__9468 (
            .O(N__42931),
            .I(\phase_controller_inst1.stoper_hc.N_318_cascade_ ));
    InMux I__9467 (
            .O(N__42928),
            .I(N__42924));
    InMux I__9466 (
            .O(N__42927),
            .I(N__42921));
    LocalMux I__9465 (
            .O(N__42924),
            .I(N__42918));
    LocalMux I__9464 (
            .O(N__42921),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    Odrv4 I__9463 (
            .O(N__42918),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__9462 (
            .O(N__42913),
            .I(N__42910));
    LocalMux I__9461 (
            .O(N__42910),
            .I(N__42906));
    InMux I__9460 (
            .O(N__42909),
            .I(N__42903));
    Odrv4 I__9459 (
            .O(N__42906),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    LocalMux I__9458 (
            .O(N__42903),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__9457 (
            .O(N__42898),
            .I(N__42895));
    LocalMux I__9456 (
            .O(N__42895),
            .I(N__42891));
    InMux I__9455 (
            .O(N__42894),
            .I(N__42888));
    Span4Mux_h I__9454 (
            .O(N__42891),
            .I(N__42885));
    LocalMux I__9453 (
            .O(N__42888),
            .I(N__42882));
    Span4Mux_v I__9452 (
            .O(N__42885),
            .I(N__42879));
    Odrv4 I__9451 (
            .O(N__42882),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    Odrv4 I__9450 (
            .O(N__42879),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    InMux I__9449 (
            .O(N__42874),
            .I(N__42871));
    LocalMux I__9448 (
            .O(N__42871),
            .I(N__42867));
    InMux I__9447 (
            .O(N__42870),
            .I(N__42863));
    Span12Mux_v I__9446 (
            .O(N__42867),
            .I(N__42860));
    InMux I__9445 (
            .O(N__42866),
            .I(N__42857));
    LocalMux I__9444 (
            .O(N__42863),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv12 I__9443 (
            .O(N__42860),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__9442 (
            .O(N__42857),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__9441 (
            .O(N__42850),
            .I(N__42847));
    LocalMux I__9440 (
            .O(N__42847),
            .I(N__42843));
    CascadeMux I__9439 (
            .O(N__42846),
            .I(N__42839));
    Span4Mux_h I__9438 (
            .O(N__42843),
            .I(N__42836));
    InMux I__9437 (
            .O(N__42842),
            .I(N__42833));
    InMux I__9436 (
            .O(N__42839),
            .I(N__42830));
    Span4Mux_h I__9435 (
            .O(N__42836),
            .I(N__42827));
    LocalMux I__9434 (
            .O(N__42833),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__9433 (
            .O(N__42830),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__9432 (
            .O(N__42827),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__9431 (
            .O(N__42820),
            .I(N__42817));
    InMux I__9430 (
            .O(N__42817),
            .I(N__42814));
    LocalMux I__9429 (
            .O(N__42814),
            .I(N__42811));
    Span4Mux_h I__9428 (
            .O(N__42811),
            .I(N__42808));
    Odrv4 I__9427 (
            .O(N__42808),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    CascadeMux I__9426 (
            .O(N__42805),
            .I(N__42802));
    InMux I__9425 (
            .O(N__42802),
            .I(N__42796));
    InMux I__9424 (
            .O(N__42801),
            .I(N__42796));
    LocalMux I__9423 (
            .O(N__42796),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    InMux I__9422 (
            .O(N__42793),
            .I(N__42790));
    LocalMux I__9421 (
            .O(N__42790),
            .I(N__42786));
    InMux I__9420 (
            .O(N__42789),
            .I(N__42783));
    Odrv4 I__9419 (
            .O(N__42786),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__9418 (
            .O(N__42783),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    CascadeMux I__9417 (
            .O(N__42778),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_ ));
    InMux I__9416 (
            .O(N__42775),
            .I(N__42770));
    InMux I__9415 (
            .O(N__42774),
            .I(N__42766));
    InMux I__9414 (
            .O(N__42773),
            .I(N__42763));
    LocalMux I__9413 (
            .O(N__42770),
            .I(N__42760));
    InMux I__9412 (
            .O(N__42769),
            .I(N__42757));
    LocalMux I__9411 (
            .O(N__42766),
            .I(N__42752));
    LocalMux I__9410 (
            .O(N__42763),
            .I(N__42752));
    Span4Mux_v I__9409 (
            .O(N__42760),
            .I(N__42749));
    LocalMux I__9408 (
            .O(N__42757),
            .I(elapsed_time_ns_1_RNIGGC6P1_0_17));
    Odrv4 I__9407 (
            .O(N__42752),
            .I(elapsed_time_ns_1_RNIGGC6P1_0_17));
    Odrv4 I__9406 (
            .O(N__42749),
            .I(elapsed_time_ns_1_RNIGGC6P1_0_17));
    CascadeMux I__9405 (
            .O(N__42742),
            .I(elapsed_time_ns_1_RNIGGC6P1_0_17_cascade_));
    CascadeMux I__9404 (
            .O(N__42739),
            .I(N__42736));
    InMux I__9403 (
            .O(N__42736),
            .I(N__42733));
    LocalMux I__9402 (
            .O(N__42733),
            .I(N__42730));
    Span4Mux_v I__9401 (
            .O(N__42730),
            .I(N__42727));
    Span4Mux_h I__9400 (
            .O(N__42727),
            .I(N__42724));
    Odrv4 I__9399 (
            .O(N__42724),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    CascadeMux I__9398 (
            .O(N__42721),
            .I(N__42718));
    InMux I__9397 (
            .O(N__42718),
            .I(N__42712));
    InMux I__9396 (
            .O(N__42717),
            .I(N__42712));
    LocalMux I__9395 (
            .O(N__42712),
            .I(N__42709));
    Span4Mux_h I__9394 (
            .O(N__42709),
            .I(N__42705));
    InMux I__9393 (
            .O(N__42708),
            .I(N__42702));
    Span4Mux_h I__9392 (
            .O(N__42705),
            .I(N__42699));
    LocalMux I__9391 (
            .O(N__42702),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__9390 (
            .O(N__42699),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__9389 (
            .O(N__42694),
            .I(N__42691));
    InMux I__9388 (
            .O(N__42691),
            .I(N__42685));
    InMux I__9387 (
            .O(N__42690),
            .I(N__42685));
    LocalMux I__9386 (
            .O(N__42685),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    InMux I__9385 (
            .O(N__42682),
            .I(N__42676));
    InMux I__9384 (
            .O(N__42681),
            .I(N__42676));
    LocalMux I__9383 (
            .O(N__42676),
            .I(N__42672));
    InMux I__9382 (
            .O(N__42675),
            .I(N__42669));
    Span12Mux_h I__9381 (
            .O(N__42672),
            .I(N__42666));
    LocalMux I__9380 (
            .O(N__42669),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv12 I__9379 (
            .O(N__42666),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__9378 (
            .O(N__42661),
            .I(N__42658));
    LocalMux I__9377 (
            .O(N__42658),
            .I(N__42655));
    Span4Mux_v I__9376 (
            .O(N__42655),
            .I(N__42652));
    Span4Mux_h I__9375 (
            .O(N__42652),
            .I(N__42649));
    Odrv4 I__9374 (
            .O(N__42649),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    InMux I__9373 (
            .O(N__42646),
            .I(N__42640));
    InMux I__9372 (
            .O(N__42645),
            .I(N__42637));
    InMux I__9371 (
            .O(N__42644),
            .I(N__42634));
    InMux I__9370 (
            .O(N__42643),
            .I(N__42631));
    LocalMux I__9369 (
            .O(N__42640),
            .I(N__42628));
    LocalMux I__9368 (
            .O(N__42637),
            .I(elapsed_time_ns_1_RNIFFC6P1_0_16));
    LocalMux I__9367 (
            .O(N__42634),
            .I(elapsed_time_ns_1_RNIFFC6P1_0_16));
    LocalMux I__9366 (
            .O(N__42631),
            .I(elapsed_time_ns_1_RNIFFC6P1_0_16));
    Odrv4 I__9365 (
            .O(N__42628),
            .I(elapsed_time_ns_1_RNIFFC6P1_0_16));
    InMux I__9364 (
            .O(N__42619),
            .I(N__42613));
    InMux I__9363 (
            .O(N__42618),
            .I(N__42613));
    LocalMux I__9362 (
            .O(N__42613),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    CascadeMux I__9361 (
            .O(N__42610),
            .I(N__42606));
    InMux I__9360 (
            .O(N__42609),
            .I(N__42601));
    InMux I__9359 (
            .O(N__42606),
            .I(N__42601));
    LocalMux I__9358 (
            .O(N__42601),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__9357 (
            .O(N__42598),
            .I(N__42595));
    LocalMux I__9356 (
            .O(N__42595),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18 ));
    CascadeMux I__9355 (
            .O(N__42592),
            .I(N__42588));
    InMux I__9354 (
            .O(N__42591),
            .I(N__42583));
    InMux I__9353 (
            .O(N__42588),
            .I(N__42583));
    LocalMux I__9352 (
            .O(N__42583),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    CascadeMux I__9351 (
            .O(N__42580),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_ ));
    InMux I__9350 (
            .O(N__42577),
            .I(N__42574));
    LocalMux I__9349 (
            .O(N__42574),
            .I(N__42570));
    InMux I__9348 (
            .O(N__42573),
            .I(N__42567));
    Odrv4 I__9347 (
            .O(N__42570),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__9346 (
            .O(N__42567),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    CascadeMux I__9345 (
            .O(N__42562),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ));
    CascadeMux I__9344 (
            .O(N__42559),
            .I(elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_));
    InMux I__9343 (
            .O(N__42556),
            .I(N__42550));
    InMux I__9342 (
            .O(N__42555),
            .I(N__42550));
    LocalMux I__9341 (
            .O(N__42550),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    InMux I__9340 (
            .O(N__42547),
            .I(N__42543));
    InMux I__9339 (
            .O(N__42546),
            .I(N__42540));
    LocalMux I__9338 (
            .O(N__42543),
            .I(N__42537));
    LocalMux I__9337 (
            .O(N__42540),
            .I(N__42534));
    Span4Mux_h I__9336 (
            .O(N__42537),
            .I(N__42531));
    Odrv4 I__9335 (
            .O(N__42534),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv4 I__9334 (
            .O(N__42531),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__9333 (
            .O(N__42526),
            .I(N__42522));
    InMux I__9332 (
            .O(N__42525),
            .I(N__42519));
    LocalMux I__9331 (
            .O(N__42522),
            .I(N__42516));
    LocalMux I__9330 (
            .O(N__42519),
            .I(N__42513));
    Span4Mux_v I__9329 (
            .O(N__42516),
            .I(N__42508));
    Span4Mux_h I__9328 (
            .O(N__42513),
            .I(N__42508));
    Odrv4 I__9327 (
            .O(N__42508),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    CascadeMux I__9326 (
            .O(N__42505),
            .I(N__42502));
    InMux I__9325 (
            .O(N__42502),
            .I(N__42499));
    LocalMux I__9324 (
            .O(N__42499),
            .I(elapsed_time_ns_1_RNIAMU8E1_0_27));
    InMux I__9323 (
            .O(N__42496),
            .I(N__42490));
    InMux I__9322 (
            .O(N__42495),
            .I(N__42490));
    LocalMux I__9321 (
            .O(N__42490),
            .I(elapsed_time_ns_1_RNI9LU8E1_0_26));
    InMux I__9320 (
            .O(N__42487),
            .I(N__42481));
    InMux I__9319 (
            .O(N__42486),
            .I(N__42481));
    LocalMux I__9318 (
            .O(N__42481),
            .I(elapsed_time_ns_1_RNIBNU8E1_0_28));
    CascadeMux I__9317 (
            .O(N__42478),
            .I(elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_));
    CascadeMux I__9316 (
            .O(N__42475),
            .I(N__42472));
    InMux I__9315 (
            .O(N__42472),
            .I(N__42468));
    InMux I__9314 (
            .O(N__42471),
            .I(N__42465));
    LocalMux I__9313 (
            .O(N__42468),
            .I(elapsed_time_ns_1_RNI8KU8E1_0_25));
    LocalMux I__9312 (
            .O(N__42465),
            .I(elapsed_time_ns_1_RNI8KU8E1_0_25));
    InMux I__9311 (
            .O(N__42460),
            .I(N__42457));
    LocalMux I__9310 (
            .O(N__42457),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15 ));
    CascadeMux I__9309 (
            .O(N__42454),
            .I(N__42451));
    InMux I__9308 (
            .O(N__42451),
            .I(N__42447));
    InMux I__9307 (
            .O(N__42450),
            .I(N__42444));
    LocalMux I__9306 (
            .O(N__42447),
            .I(elapsed_time_ns_1_RNI5HU8E1_0_22));
    LocalMux I__9305 (
            .O(N__42444),
            .I(elapsed_time_ns_1_RNI5HU8E1_0_22));
    CascadeMux I__9304 (
            .O(N__42439),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15_cascade_ ));
    CascadeMux I__9303 (
            .O(N__42436),
            .I(N__42433));
    InMux I__9302 (
            .O(N__42433),
            .I(N__42429));
    InMux I__9301 (
            .O(N__42432),
            .I(N__42426));
    LocalMux I__9300 (
            .O(N__42429),
            .I(elapsed_time_ns_1_RNI7JU8E1_0_24));
    LocalMux I__9299 (
            .O(N__42426),
            .I(elapsed_time_ns_1_RNI7JU8E1_0_24));
    CascadeMux I__9298 (
            .O(N__42421),
            .I(N__42418));
    InMux I__9297 (
            .O(N__42418),
            .I(N__42414));
    InMux I__9296 (
            .O(N__42417),
            .I(N__42411));
    LocalMux I__9295 (
            .O(N__42414),
            .I(elapsed_time_ns_1_RNI6IU8E1_0_23));
    LocalMux I__9294 (
            .O(N__42411),
            .I(elapsed_time_ns_1_RNI6IU8E1_0_23));
    InMux I__9293 (
            .O(N__42406),
            .I(N__42403));
    LocalMux I__9292 (
            .O(N__42403),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15 ));
    InMux I__9291 (
            .O(N__42400),
            .I(N__42396));
    InMux I__9290 (
            .O(N__42399),
            .I(N__42393));
    LocalMux I__9289 (
            .O(N__42396),
            .I(N__42390));
    LocalMux I__9288 (
            .O(N__42393),
            .I(N__42387));
    Odrv4 I__9287 (
            .O(N__42390),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__9286 (
            .O(N__42387),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__9285 (
            .O(N__42382),
            .I(N__42379));
    LocalMux I__9284 (
            .O(N__42379),
            .I(N__42375));
    InMux I__9283 (
            .O(N__42378),
            .I(N__42372));
    Odrv4 I__9282 (
            .O(N__42375),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__9281 (
            .O(N__42372),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__9280 (
            .O(N__42367),
            .I(N__42364));
    LocalMux I__9279 (
            .O(N__42364),
            .I(N__42360));
    InMux I__9278 (
            .O(N__42363),
            .I(N__42357));
    Odrv4 I__9277 (
            .O(N__42360),
            .I(\delay_measurement_inst.delay_hc_timer.N_369 ));
    LocalMux I__9276 (
            .O(N__42357),
            .I(\delay_measurement_inst.delay_hc_timer.N_369 ));
    CascadeMux I__9275 (
            .O(N__42352),
            .I(\delay_measurement_inst.delay_hc_timer.N_344_i_cascade_ ));
    CascadeMux I__9274 (
            .O(N__42349),
            .I(elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_));
    InMux I__9273 (
            .O(N__42346),
            .I(N__42340));
    InMux I__9272 (
            .O(N__42345),
            .I(N__42340));
    LocalMux I__9271 (
            .O(N__42340),
            .I(N__42337));
    Span4Mux_h I__9270 (
            .O(N__42337),
            .I(N__42334));
    Odrv4 I__9269 (
            .O(N__42334),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__9268 (
            .O(N__42331),
            .I(N__42328));
    LocalMux I__9267 (
            .O(N__42328),
            .I(N__42324));
    InMux I__9266 (
            .O(N__42327),
            .I(N__42321));
    Span4Mux_h I__9265 (
            .O(N__42324),
            .I(N__42318));
    LocalMux I__9264 (
            .O(N__42321),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__9263 (
            .O(N__42318),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    CascadeMux I__9262 (
            .O(N__42313),
            .I(N__42310));
    InMux I__9261 (
            .O(N__42310),
            .I(N__42307));
    LocalMux I__9260 (
            .O(N__42307),
            .I(N__42303));
    InMux I__9259 (
            .O(N__42306),
            .I(N__42299));
    Span4Mux_h I__9258 (
            .O(N__42303),
            .I(N__42296));
    InMux I__9257 (
            .O(N__42302),
            .I(N__42293));
    LocalMux I__9256 (
            .O(N__42299),
            .I(elapsed_time_ns_1_RNIMHKEE1_0_5));
    Odrv4 I__9255 (
            .O(N__42296),
            .I(elapsed_time_ns_1_RNIMHKEE1_0_5));
    LocalMux I__9254 (
            .O(N__42293),
            .I(elapsed_time_ns_1_RNIMHKEE1_0_5));
    InMux I__9253 (
            .O(N__42286),
            .I(N__42276));
    CascadeMux I__9252 (
            .O(N__42285),
            .I(N__42273));
    InMux I__9251 (
            .O(N__42284),
            .I(N__42268));
    InMux I__9250 (
            .O(N__42283),
            .I(N__42256));
    InMux I__9249 (
            .O(N__42282),
            .I(N__42256));
    InMux I__9248 (
            .O(N__42281),
            .I(N__42256));
    InMux I__9247 (
            .O(N__42280),
            .I(N__42256));
    InMux I__9246 (
            .O(N__42279),
            .I(N__42256));
    LocalMux I__9245 (
            .O(N__42276),
            .I(N__42253));
    InMux I__9244 (
            .O(N__42273),
            .I(N__42248));
    InMux I__9243 (
            .O(N__42272),
            .I(N__42248));
    InMux I__9242 (
            .O(N__42271),
            .I(N__42245));
    LocalMux I__9241 (
            .O(N__42268),
            .I(N__42242));
    InMux I__9240 (
            .O(N__42267),
            .I(N__42239));
    LocalMux I__9239 (
            .O(N__42256),
            .I(N__42228));
    Span4Mux_h I__9238 (
            .O(N__42253),
            .I(N__42228));
    LocalMux I__9237 (
            .O(N__42248),
            .I(N__42228));
    LocalMux I__9236 (
            .O(N__42245),
            .I(N__42228));
    Span4Mux_h I__9235 (
            .O(N__42242),
            .I(N__42228));
    LocalMux I__9234 (
            .O(N__42239),
            .I(\phase_controller_inst1.stoper_hc.N_330 ));
    Odrv4 I__9233 (
            .O(N__42228),
            .I(\phase_controller_inst1.stoper_hc.N_330 ));
    CascadeMux I__9232 (
            .O(N__42223),
            .I(elapsed_time_ns_1_RNIMHKEE1_0_5_cascade_));
    CascadeMux I__9231 (
            .O(N__42220),
            .I(N__42217));
    InMux I__9230 (
            .O(N__42217),
            .I(N__42209));
    InMux I__9229 (
            .O(N__42216),
            .I(N__42206));
    CascadeMux I__9228 (
            .O(N__42215),
            .I(N__42197));
    CascadeMux I__9227 (
            .O(N__42214),
            .I(N__42194));
    InMux I__9226 (
            .O(N__42213),
            .I(N__42189));
    InMux I__9225 (
            .O(N__42212),
            .I(N__42186));
    LocalMux I__9224 (
            .O(N__42209),
            .I(N__42181));
    LocalMux I__9223 (
            .O(N__42206),
            .I(N__42181));
    InMux I__9222 (
            .O(N__42205),
            .I(N__42178));
    InMux I__9221 (
            .O(N__42204),
            .I(N__42173));
    InMux I__9220 (
            .O(N__42203),
            .I(N__42173));
    InMux I__9219 (
            .O(N__42202),
            .I(N__42162));
    InMux I__9218 (
            .O(N__42201),
            .I(N__42162));
    InMux I__9217 (
            .O(N__42200),
            .I(N__42162));
    InMux I__9216 (
            .O(N__42197),
            .I(N__42162));
    InMux I__9215 (
            .O(N__42194),
            .I(N__42162));
    InMux I__9214 (
            .O(N__42193),
            .I(N__42157));
    InMux I__9213 (
            .O(N__42192),
            .I(N__42157));
    LocalMux I__9212 (
            .O(N__42189),
            .I(N__42154));
    LocalMux I__9211 (
            .O(N__42186),
            .I(N__42149));
    Span4Mux_h I__9210 (
            .O(N__42181),
            .I(N__42149));
    LocalMux I__9209 (
            .O(N__42178),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    LocalMux I__9208 (
            .O(N__42173),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    LocalMux I__9207 (
            .O(N__42162),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    LocalMux I__9206 (
            .O(N__42157),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    Odrv4 I__9205 (
            .O(N__42154),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    Odrv4 I__9204 (
            .O(N__42149),
            .I(\phase_controller_inst1.stoper_hc.N_328 ));
    InMux I__9203 (
            .O(N__42136),
            .I(N__42132));
    InMux I__9202 (
            .O(N__42135),
            .I(N__42129));
    LocalMux I__9201 (
            .O(N__42132),
            .I(N__42124));
    LocalMux I__9200 (
            .O(N__42129),
            .I(N__42124));
    Span4Mux_v I__9199 (
            .O(N__42124),
            .I(N__42121));
    Odrv4 I__9198 (
            .O(N__42121),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__9197 (
            .O(N__42118),
            .I(N__42114));
    InMux I__9196 (
            .O(N__42117),
            .I(N__42111));
    LocalMux I__9195 (
            .O(N__42114),
            .I(N__42106));
    LocalMux I__9194 (
            .O(N__42111),
            .I(N__42106));
    Odrv4 I__9193 (
            .O(N__42106),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    CascadeMux I__9192 (
            .O(N__42103),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19_cascade_ ));
    CascadeMux I__9191 (
            .O(N__42100),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_ ));
    CascadeMux I__9190 (
            .O(N__42097),
            .I(elapsed_time_ns_1_RNI4FT8E1_0_12_cascade_));
    InMux I__9189 (
            .O(N__42094),
            .I(N__42091));
    LocalMux I__9188 (
            .O(N__42091),
            .I(N__42088));
    Span4Mux_h I__9187 (
            .O(N__42088),
            .I(N__42085));
    Odrv4 I__9186 (
            .O(N__42085),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15 ));
    InMux I__9185 (
            .O(N__42082),
            .I(N__42079));
    LocalMux I__9184 (
            .O(N__42079),
            .I(N__42076));
    Span4Mux_h I__9183 (
            .O(N__42076),
            .I(N__42073));
    Odrv4 I__9182 (
            .O(N__42073),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14 ));
    CascadeMux I__9181 (
            .O(N__42070),
            .I(N__42067));
    InMux I__9180 (
            .O(N__42067),
            .I(N__42064));
    LocalMux I__9179 (
            .O(N__42064),
            .I(N__42061));
    Span4Mux_h I__9178 (
            .O(N__42061),
            .I(N__42058));
    Odrv4 I__9177 (
            .O(N__42058),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20 ));
    CascadeMux I__9176 (
            .O(N__42055),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_ ));
    CascadeMux I__9175 (
            .O(N__42052),
            .I(\delay_measurement_inst.delay_hc_timer.N_369_cascade_ ));
    CascadeMux I__9174 (
            .O(N__42049),
            .I(\delay_measurement_inst.delay_hc_timer.N_367_clk_cascade_ ));
    InMux I__9173 (
            .O(N__42046),
            .I(N__42042));
    InMux I__9172 (
            .O(N__42045),
            .I(N__42039));
    LocalMux I__9171 (
            .O(N__42042),
            .I(elapsed_time_ns_1_RNI3FU8E1_0_20));
    LocalMux I__9170 (
            .O(N__42039),
            .I(elapsed_time_ns_1_RNI3FU8E1_0_20));
    InMux I__9169 (
            .O(N__42034),
            .I(N__42030));
    InMux I__9168 (
            .O(N__42033),
            .I(N__42027));
    LocalMux I__9167 (
            .O(N__42030),
            .I(N__42024));
    LocalMux I__9166 (
            .O(N__42027),
            .I(N__42021));
    Odrv12 I__9165 (
            .O(N__42024),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv4 I__9164 (
            .O(N__42021),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    CascadeMux I__9163 (
            .O(N__42016),
            .I(N__42012));
    InMux I__9162 (
            .O(N__42015),
            .I(N__42009));
    InMux I__9161 (
            .O(N__42012),
            .I(N__42006));
    LocalMux I__9160 (
            .O(N__42009),
            .I(N__42003));
    LocalMux I__9159 (
            .O(N__42006),
            .I(N__42000));
    Span4Mux_v I__9158 (
            .O(N__42003),
            .I(N__41997));
    Span4Mux_h I__9157 (
            .O(N__42000),
            .I(N__41994));
    Odrv4 I__9156 (
            .O(N__41997),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    Odrv4 I__9155 (
            .O(N__41994),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    CascadeMux I__9154 (
            .O(N__41989),
            .I(N__41986));
    InMux I__9153 (
            .O(N__41986),
            .I(N__41983));
    LocalMux I__9152 (
            .O(N__41983),
            .I(N__41980));
    Span4Mux_h I__9151 (
            .O(N__41980),
            .I(N__41977));
    Odrv4 I__9150 (
            .O(N__41977),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    InMux I__9149 (
            .O(N__41974),
            .I(N__41971));
    LocalMux I__9148 (
            .O(N__41971),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    InMux I__9147 (
            .O(N__41968),
            .I(N__41964));
    InMux I__9146 (
            .O(N__41967),
            .I(N__41960));
    LocalMux I__9145 (
            .O(N__41964),
            .I(N__41957));
    InMux I__9144 (
            .O(N__41963),
            .I(N__41952));
    LocalMux I__9143 (
            .O(N__41960),
            .I(N__41949));
    Span4Mux_h I__9142 (
            .O(N__41957),
            .I(N__41946));
    InMux I__9141 (
            .O(N__41956),
            .I(N__41941));
    InMux I__9140 (
            .O(N__41955),
            .I(N__41941));
    LocalMux I__9139 (
            .O(N__41952),
            .I(elapsed_time_ns_1_RNI8765M1_0_16));
    Odrv12 I__9138 (
            .O(N__41949),
            .I(elapsed_time_ns_1_RNI8765M1_0_16));
    Odrv4 I__9137 (
            .O(N__41946),
            .I(elapsed_time_ns_1_RNI8765M1_0_16));
    LocalMux I__9136 (
            .O(N__41941),
            .I(elapsed_time_ns_1_RNI8765M1_0_16));
    InMux I__9135 (
            .O(N__41932),
            .I(N__41926));
    InMux I__9134 (
            .O(N__41931),
            .I(N__41926));
    LocalMux I__9133 (
            .O(N__41926),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__9132 (
            .O(N__41923),
            .I(N__41919));
    InMux I__9131 (
            .O(N__41922),
            .I(N__41915));
    LocalMux I__9130 (
            .O(N__41919),
            .I(N__41912));
    CascadeMux I__9129 (
            .O(N__41918),
            .I(N__41908));
    LocalMux I__9128 (
            .O(N__41915),
            .I(N__41905));
    Span4Mux_h I__9127 (
            .O(N__41912),
            .I(N__41902));
    InMux I__9126 (
            .O(N__41911),
            .I(N__41899));
    InMux I__9125 (
            .O(N__41908),
            .I(N__41896));
    Odrv4 I__9124 (
            .O(N__41905),
            .I(elapsed_time_ns_1_RNI9865M1_0_17));
    Odrv4 I__9123 (
            .O(N__41902),
            .I(elapsed_time_ns_1_RNI9865M1_0_17));
    LocalMux I__9122 (
            .O(N__41899),
            .I(elapsed_time_ns_1_RNI9865M1_0_17));
    LocalMux I__9121 (
            .O(N__41896),
            .I(elapsed_time_ns_1_RNI9865M1_0_17));
    CascadeMux I__9120 (
            .O(N__41887),
            .I(N__41884));
    InMux I__9119 (
            .O(N__41884),
            .I(N__41878));
    InMux I__9118 (
            .O(N__41883),
            .I(N__41878));
    LocalMux I__9117 (
            .O(N__41878),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__9116 (
            .O(N__41875),
            .I(N__41869));
    InMux I__9115 (
            .O(N__41874),
            .I(N__41869));
    LocalMux I__9114 (
            .O(N__41869),
            .I(N__41865));
    InMux I__9113 (
            .O(N__41868),
            .I(N__41862));
    Span4Mux_h I__9112 (
            .O(N__41865),
            .I(N__41857));
    LocalMux I__9111 (
            .O(N__41862),
            .I(N__41854));
    InMux I__9110 (
            .O(N__41861),
            .I(N__41851));
    InMux I__9109 (
            .O(N__41860),
            .I(N__41848));
    Odrv4 I__9108 (
            .O(N__41857),
            .I(elapsed_time_ns_1_RNIBA65M1_0_19));
    Odrv4 I__9107 (
            .O(N__41854),
            .I(elapsed_time_ns_1_RNIBA65M1_0_19));
    LocalMux I__9106 (
            .O(N__41851),
            .I(elapsed_time_ns_1_RNIBA65M1_0_19));
    LocalMux I__9105 (
            .O(N__41848),
            .I(elapsed_time_ns_1_RNIBA65M1_0_19));
    CascadeMux I__9104 (
            .O(N__41839),
            .I(N__41836));
    InMux I__9103 (
            .O(N__41836),
            .I(N__41833));
    LocalMux I__9102 (
            .O(N__41833),
            .I(N__41830));
    Odrv4 I__9101 (
            .O(N__41830),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    CascadeMux I__9100 (
            .O(N__41827),
            .I(N__41824));
    InMux I__9099 (
            .O(N__41824),
            .I(N__41818));
    InMux I__9098 (
            .O(N__41823),
            .I(N__41818));
    LocalMux I__9097 (
            .O(N__41818),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__9096 (
            .O(N__41815),
            .I(N__41812));
    LocalMux I__9095 (
            .O(N__41812),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__9094 (
            .O(N__41809),
            .I(N__41787));
    InMux I__9093 (
            .O(N__41808),
            .I(N__41787));
    InMux I__9092 (
            .O(N__41807),
            .I(N__41787));
    InMux I__9091 (
            .O(N__41806),
            .I(N__41787));
    InMux I__9090 (
            .O(N__41805),
            .I(N__41787));
    InMux I__9089 (
            .O(N__41804),
            .I(N__41782));
    InMux I__9088 (
            .O(N__41803),
            .I(N__41782));
    CascadeMux I__9087 (
            .O(N__41802),
            .I(N__41765));
    InMux I__9086 (
            .O(N__41801),
            .I(N__41752));
    InMux I__9085 (
            .O(N__41800),
            .I(N__41752));
    InMux I__9084 (
            .O(N__41799),
            .I(N__41752));
    InMux I__9083 (
            .O(N__41798),
            .I(N__41752));
    LocalMux I__9082 (
            .O(N__41787),
            .I(N__41746));
    LocalMux I__9081 (
            .O(N__41782),
            .I(N__41743));
    InMux I__9080 (
            .O(N__41781),
            .I(N__41732));
    InMux I__9079 (
            .O(N__41780),
            .I(N__41732));
    InMux I__9078 (
            .O(N__41779),
            .I(N__41732));
    InMux I__9077 (
            .O(N__41778),
            .I(N__41732));
    InMux I__9076 (
            .O(N__41777),
            .I(N__41732));
    InMux I__9075 (
            .O(N__41776),
            .I(N__41719));
    InMux I__9074 (
            .O(N__41775),
            .I(N__41719));
    InMux I__9073 (
            .O(N__41774),
            .I(N__41719));
    InMux I__9072 (
            .O(N__41773),
            .I(N__41719));
    InMux I__9071 (
            .O(N__41772),
            .I(N__41719));
    InMux I__9070 (
            .O(N__41771),
            .I(N__41719));
    InMux I__9069 (
            .O(N__41770),
            .I(N__41716));
    InMux I__9068 (
            .O(N__41769),
            .I(N__41707));
    InMux I__9067 (
            .O(N__41768),
            .I(N__41707));
    InMux I__9066 (
            .O(N__41765),
            .I(N__41707));
    InMux I__9065 (
            .O(N__41764),
            .I(N__41707));
    InMux I__9064 (
            .O(N__41763),
            .I(N__41700));
    InMux I__9063 (
            .O(N__41762),
            .I(N__41700));
    InMux I__9062 (
            .O(N__41761),
            .I(N__41700));
    LocalMux I__9061 (
            .O(N__41752),
            .I(N__41695));
    InMux I__9060 (
            .O(N__41751),
            .I(N__41688));
    InMux I__9059 (
            .O(N__41750),
            .I(N__41688));
    InMux I__9058 (
            .O(N__41749),
            .I(N__41688));
    Span4Mux_v I__9057 (
            .O(N__41746),
            .I(N__41681));
    Span4Mux_v I__9056 (
            .O(N__41743),
            .I(N__41681));
    LocalMux I__9055 (
            .O(N__41732),
            .I(N__41681));
    LocalMux I__9054 (
            .O(N__41719),
            .I(N__41672));
    LocalMux I__9053 (
            .O(N__41716),
            .I(N__41672));
    LocalMux I__9052 (
            .O(N__41707),
            .I(N__41672));
    LocalMux I__9051 (
            .O(N__41700),
            .I(N__41672));
    InMux I__9050 (
            .O(N__41699),
            .I(N__41667));
    InMux I__9049 (
            .O(N__41698),
            .I(N__41667));
    Odrv4 I__9048 (
            .O(N__41695),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__9047 (
            .O(N__41688),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__9046 (
            .O(N__41681),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    Odrv4 I__9045 (
            .O(N__41672),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    LocalMux I__9044 (
            .O(N__41667),
            .I(elapsed_time_ns_1_RNISCJF91_0_31));
    CascadeMux I__9043 (
            .O(N__41656),
            .I(N__41652));
    CascadeMux I__9042 (
            .O(N__41655),
            .I(N__41649));
    InMux I__9041 (
            .O(N__41652),
            .I(N__41638));
    InMux I__9040 (
            .O(N__41649),
            .I(N__41638));
    InMux I__9039 (
            .O(N__41648),
            .I(N__41638));
    InMux I__9038 (
            .O(N__41647),
            .I(N__41638));
    LocalMux I__9037 (
            .O(N__41638),
            .I(N__41618));
    InMux I__9036 (
            .O(N__41637),
            .I(N__41607));
    InMux I__9035 (
            .O(N__41636),
            .I(N__41607));
    InMux I__9034 (
            .O(N__41635),
            .I(N__41607));
    InMux I__9033 (
            .O(N__41634),
            .I(N__41607));
    InMux I__9032 (
            .O(N__41633),
            .I(N__41607));
    CascadeMux I__9031 (
            .O(N__41632),
            .I(N__41604));
    CascadeMux I__9030 (
            .O(N__41631),
            .I(N__41601));
    CascadeMux I__9029 (
            .O(N__41630),
            .I(N__41597));
    InMux I__9028 (
            .O(N__41629),
            .I(N__41586));
    InMux I__9027 (
            .O(N__41628),
            .I(N__41586));
    InMux I__9026 (
            .O(N__41627),
            .I(N__41586));
    InMux I__9025 (
            .O(N__41626),
            .I(N__41583));
    InMux I__9024 (
            .O(N__41625),
            .I(N__41578));
    InMux I__9023 (
            .O(N__41624),
            .I(N__41578));
    CascadeMux I__9022 (
            .O(N__41623),
            .I(N__41575));
    CascadeMux I__9021 (
            .O(N__41622),
            .I(N__41572));
    CascadeMux I__9020 (
            .O(N__41621),
            .I(N__41569));
    Span4Mux_h I__9019 (
            .O(N__41618),
            .I(N__41565));
    LocalMux I__9018 (
            .O(N__41607),
            .I(N__41562));
    InMux I__9017 (
            .O(N__41604),
            .I(N__41555));
    InMux I__9016 (
            .O(N__41601),
            .I(N__41555));
    InMux I__9015 (
            .O(N__41600),
            .I(N__41555));
    InMux I__9014 (
            .O(N__41597),
            .I(N__41546));
    InMux I__9013 (
            .O(N__41596),
            .I(N__41546));
    InMux I__9012 (
            .O(N__41595),
            .I(N__41546));
    InMux I__9011 (
            .O(N__41594),
            .I(N__41546));
    InMux I__9010 (
            .O(N__41593),
            .I(N__41543));
    LocalMux I__9009 (
            .O(N__41586),
            .I(N__41538));
    LocalMux I__9008 (
            .O(N__41583),
            .I(N__41538));
    LocalMux I__9007 (
            .O(N__41578),
            .I(N__41535));
    InMux I__9006 (
            .O(N__41575),
            .I(N__41526));
    InMux I__9005 (
            .O(N__41572),
            .I(N__41526));
    InMux I__9004 (
            .O(N__41569),
            .I(N__41526));
    InMux I__9003 (
            .O(N__41568),
            .I(N__41526));
    Span4Mux_v I__9002 (
            .O(N__41565),
            .I(N__41521));
    Span4Mux_h I__9001 (
            .O(N__41562),
            .I(N__41521));
    LocalMux I__9000 (
            .O(N__41555),
            .I(N__41510));
    LocalMux I__8999 (
            .O(N__41546),
            .I(N__41510));
    LocalMux I__8998 (
            .O(N__41543),
            .I(N__41510));
    Span4Mux_v I__8997 (
            .O(N__41538),
            .I(N__41510));
    Span4Mux_h I__8996 (
            .O(N__41535),
            .I(N__41510));
    LocalMux I__8995 (
            .O(N__41526),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv4 I__8994 (
            .O(N__41521),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    Odrv4 I__8993 (
            .O(N__41510),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ));
    InMux I__8992 (
            .O(N__41503),
            .I(N__41499));
    InMux I__8991 (
            .O(N__41502),
            .I(N__41495));
    LocalMux I__8990 (
            .O(N__41499),
            .I(N__41492));
    CascadeMux I__8989 (
            .O(N__41498),
            .I(N__41489));
    LocalMux I__8988 (
            .O(N__41495),
            .I(N__41485));
    Span4Mux_h I__8987 (
            .O(N__41492),
            .I(N__41482));
    InMux I__8986 (
            .O(N__41489),
            .I(N__41479));
    InMux I__8985 (
            .O(N__41488),
            .I(N__41476));
    Odrv4 I__8984 (
            .O(N__41485),
            .I(elapsed_time_ns_1_RNIA965M1_0_18));
    Odrv4 I__8983 (
            .O(N__41482),
            .I(elapsed_time_ns_1_RNIA965M1_0_18));
    LocalMux I__8982 (
            .O(N__41479),
            .I(elapsed_time_ns_1_RNIA965M1_0_18));
    LocalMux I__8981 (
            .O(N__41476),
            .I(elapsed_time_ns_1_RNIA965M1_0_18));
    InMux I__8980 (
            .O(N__41467),
            .I(N__41461));
    InMux I__8979 (
            .O(N__41466),
            .I(N__41461));
    LocalMux I__8978 (
            .O(N__41461),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__8977 (
            .O(N__41458),
            .I(N__41455));
    LocalMux I__8976 (
            .O(N__41455),
            .I(N__41452));
    Odrv4 I__8975 (
            .O(N__41452),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14 ));
    CascadeMux I__8974 (
            .O(N__41449),
            .I(N__41445));
    InMux I__8973 (
            .O(N__41448),
            .I(N__41440));
    InMux I__8972 (
            .O(N__41445),
            .I(N__41437));
    InMux I__8971 (
            .O(N__41444),
            .I(N__41434));
    InMux I__8970 (
            .O(N__41443),
            .I(N__41429));
    LocalMux I__8969 (
            .O(N__41440),
            .I(N__41426));
    LocalMux I__8968 (
            .O(N__41437),
            .I(N__41421));
    LocalMux I__8967 (
            .O(N__41434),
            .I(N__41421));
    InMux I__8966 (
            .O(N__41433),
            .I(N__41418));
    InMux I__8965 (
            .O(N__41432),
            .I(N__41415));
    LocalMux I__8964 (
            .O(N__41429),
            .I(N__41412));
    Span4Mux_h I__8963 (
            .O(N__41426),
            .I(N__41409));
    Span4Mux_v I__8962 (
            .O(N__41421),
            .I(N__41402));
    LocalMux I__8961 (
            .O(N__41418),
            .I(N__41402));
    LocalMux I__8960 (
            .O(N__41415),
            .I(N__41402));
    Odrv12 I__8959 (
            .O(N__41412),
            .I(elapsed_time_ns_1_RNI6565M1_0_14));
    Odrv4 I__8958 (
            .O(N__41409),
            .I(elapsed_time_ns_1_RNI6565M1_0_14));
    Odrv4 I__8957 (
            .O(N__41402),
            .I(elapsed_time_ns_1_RNI6565M1_0_14));
    InMux I__8956 (
            .O(N__41395),
            .I(N__41392));
    LocalMux I__8955 (
            .O(N__41392),
            .I(N__41388));
    InMux I__8954 (
            .O(N__41391),
            .I(N__41385));
    Odrv12 I__8953 (
            .O(N__41388),
            .I(\delay_measurement_inst.delay_tr_timer.N_395 ));
    LocalMux I__8952 (
            .O(N__41385),
            .I(\delay_measurement_inst.delay_tr_timer.N_395 ));
    InMux I__8951 (
            .O(N__41380),
            .I(N__41377));
    LocalMux I__8950 (
            .O(N__41377),
            .I(N__41373));
    InMux I__8949 (
            .O(N__41376),
            .I(N__41370));
    Odrv4 I__8948 (
            .O(N__41373),
            .I(\delay_measurement_inst.delay_tr_timer.N_375 ));
    LocalMux I__8947 (
            .O(N__41370),
            .I(\delay_measurement_inst.delay_tr_timer.N_375 ));
    InMux I__8946 (
            .O(N__41365),
            .I(N__41355));
    InMux I__8945 (
            .O(N__41364),
            .I(N__41348));
    InMux I__8944 (
            .O(N__41363),
            .I(N__41348));
    InMux I__8943 (
            .O(N__41362),
            .I(N__41348));
    InMux I__8942 (
            .O(N__41361),
            .I(N__41339));
    InMux I__8941 (
            .O(N__41360),
            .I(N__41339));
    InMux I__8940 (
            .O(N__41359),
            .I(N__41339));
    InMux I__8939 (
            .O(N__41358),
            .I(N__41339));
    LocalMux I__8938 (
            .O(N__41355),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    LocalMux I__8937 (
            .O(N__41348),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    LocalMux I__8936 (
            .O(N__41339),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ));
    InMux I__8935 (
            .O(N__41332),
            .I(N__41329));
    LocalMux I__8934 (
            .O(N__41329),
            .I(N__41326));
    Odrv4 I__8933 (
            .O(N__41326),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ));
    CascadeMux I__8932 (
            .O(N__41323),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ));
    InMux I__8931 (
            .O(N__41320),
            .I(N__41312));
    InMux I__8930 (
            .O(N__41319),
            .I(N__41312));
    InMux I__8929 (
            .O(N__41318),
            .I(N__41307));
    InMux I__8928 (
            .O(N__41317),
            .I(N__41304));
    LocalMux I__8927 (
            .O(N__41312),
            .I(N__41301));
    InMux I__8926 (
            .O(N__41311),
            .I(N__41296));
    InMux I__8925 (
            .O(N__41310),
            .I(N__41296));
    LocalMux I__8924 (
            .O(N__41307),
            .I(N__41291));
    LocalMux I__8923 (
            .O(N__41304),
            .I(N__41291));
    Span4Mux_v I__8922 (
            .O(N__41301),
            .I(N__41286));
    LocalMux I__8921 (
            .O(N__41296),
            .I(N__41286));
    Odrv4 I__8920 (
            .O(N__41291),
            .I(elapsed_time_ns_1_RNIQENQL1_0_9));
    Odrv4 I__8919 (
            .O(N__41286),
            .I(elapsed_time_ns_1_RNIQENQL1_0_9));
    CascadeMux I__8918 (
            .O(N__41281),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_ ));
    InMux I__8917 (
            .O(N__41278),
            .I(N__41275));
    LocalMux I__8916 (
            .O(N__41275),
            .I(N__41271));
    InMux I__8915 (
            .O(N__41274),
            .I(N__41268));
    Odrv12 I__8914 (
            .O(N__41271),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    LocalMux I__8913 (
            .O(N__41268),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    InMux I__8912 (
            .O(N__41263),
            .I(N__41256));
    InMux I__8911 (
            .O(N__41262),
            .I(N__41256));
    InMux I__8910 (
            .O(N__41261),
            .I(N__41253));
    LocalMux I__8909 (
            .O(N__41256),
            .I(N__41250));
    LocalMux I__8908 (
            .O(N__41253),
            .I(N__41247));
    Span4Mux_h I__8907 (
            .O(N__41250),
            .I(N__41243));
    Span4Mux_v I__8906 (
            .O(N__41247),
            .I(N__41240));
    InMux I__8905 (
            .O(N__41246),
            .I(N__41237));
    Span4Mux_v I__8904 (
            .O(N__41243),
            .I(N__41234));
    Odrv4 I__8903 (
            .O(N__41240),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__8902 (
            .O(N__41237),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv4 I__8901 (
            .O(N__41234),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    CascadeMux I__8900 (
            .O(N__41227),
            .I(N__41224));
    InMux I__8899 (
            .O(N__41224),
            .I(N__41219));
    InMux I__8898 (
            .O(N__41223),
            .I(N__41214));
    InMux I__8897 (
            .O(N__41222),
            .I(N__41214));
    LocalMux I__8896 (
            .O(N__41219),
            .I(N__41211));
    LocalMux I__8895 (
            .O(N__41214),
            .I(N__41208));
    Span12Mux_h I__8894 (
            .O(N__41211),
            .I(N__41205));
    Span12Mux_v I__8893 (
            .O(N__41208),
            .I(N__41200));
    Span12Mux_v I__8892 (
            .O(N__41205),
            .I(N__41200));
    Odrv12 I__8891 (
            .O(N__41200),
            .I(il_max_comp2_D2));
    InMux I__8890 (
            .O(N__41197),
            .I(N__41194));
    LocalMux I__8889 (
            .O(N__41194),
            .I(N__41191));
    Span4Mux_h I__8888 (
            .O(N__41191),
            .I(N__41186));
    InMux I__8887 (
            .O(N__41190),
            .I(N__41181));
    InMux I__8886 (
            .O(N__41189),
            .I(N__41181));
    Odrv4 I__8885 (
            .O(N__41186),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__8884 (
            .O(N__41181),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    CascadeMux I__8883 (
            .O(N__41176),
            .I(\delay_measurement_inst.delay_tr_timer.N_353_cascade_ ));
    InMux I__8882 (
            .O(N__41173),
            .I(N__41170));
    LocalMux I__8881 (
            .O(N__41170),
            .I(N__41165));
    InMux I__8880 (
            .O(N__41169),
            .I(N__41160));
    InMux I__8879 (
            .O(N__41168),
            .I(N__41160));
    Odrv4 I__8878 (
            .O(N__41165),
            .I(\delay_measurement_inst.delay_tr_timer.N_382 ));
    LocalMux I__8877 (
            .O(N__41160),
            .I(\delay_measurement_inst.delay_tr_timer.N_382 ));
    InMux I__8876 (
            .O(N__41155),
            .I(N__41152));
    LocalMux I__8875 (
            .O(N__41152),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16 ));
    InMux I__8874 (
            .O(N__41149),
            .I(N__41146));
    LocalMux I__8873 (
            .O(N__41146),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ));
    CascadeMux I__8872 (
            .O(N__41143),
            .I(N__41140));
    InMux I__8871 (
            .O(N__41140),
            .I(N__41135));
    CascadeMux I__8870 (
            .O(N__41139),
            .I(N__41132));
    InMux I__8869 (
            .O(N__41138),
            .I(N__41129));
    LocalMux I__8868 (
            .O(N__41135),
            .I(N__41126));
    InMux I__8867 (
            .O(N__41132),
            .I(N__41122));
    LocalMux I__8866 (
            .O(N__41129),
            .I(N__41117));
    Span4Mux_h I__8865 (
            .O(N__41126),
            .I(N__41117));
    InMux I__8864 (
            .O(N__41125),
            .I(N__41114));
    LocalMux I__8863 (
            .O(N__41122),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    Odrv4 I__8862 (
            .O(N__41117),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    LocalMux I__8861 (
            .O(N__41114),
            .I(elapsed_time_ns_1_RNIDH2591_0_5));
    CascadeMux I__8860 (
            .O(N__41107),
            .I(elapsed_time_ns_1_RNIA965M1_0_18_cascade_));
    CascadeMux I__8859 (
            .O(N__41104),
            .I(N__41101));
    InMux I__8858 (
            .O(N__41101),
            .I(N__41097));
    InMux I__8857 (
            .O(N__41100),
            .I(N__41093));
    LocalMux I__8856 (
            .O(N__41097),
            .I(N__41090));
    InMux I__8855 (
            .O(N__41096),
            .I(N__41086));
    LocalMux I__8854 (
            .O(N__41093),
            .I(N__41083));
    Span4Mux_v I__8853 (
            .O(N__41090),
            .I(N__41080));
    InMux I__8852 (
            .O(N__41089),
            .I(N__41077));
    LocalMux I__8851 (
            .O(N__41086),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    Odrv4 I__8850 (
            .O(N__41083),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    Odrv4 I__8849 (
            .O(N__41080),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    LocalMux I__8848 (
            .O(N__41077),
            .I(elapsed_time_ns_1_RNICG2591_0_4));
    InMux I__8847 (
            .O(N__41068),
            .I(N__41065));
    LocalMux I__8846 (
            .O(N__41065),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2 ));
    CascadeMux I__8845 (
            .O(N__41062),
            .I(N__41057));
    CascadeMux I__8844 (
            .O(N__41061),
            .I(N__41051));
    CascadeMux I__8843 (
            .O(N__41060),
            .I(N__41046));
    InMux I__8842 (
            .O(N__41057),
            .I(N__41036));
    InMux I__8841 (
            .O(N__41056),
            .I(N__41026));
    InMux I__8840 (
            .O(N__41055),
            .I(N__41019));
    InMux I__8839 (
            .O(N__41054),
            .I(N__41014));
    InMux I__8838 (
            .O(N__41051),
            .I(N__41014));
    CascadeMux I__8837 (
            .O(N__41050),
            .I(N__41011));
    CascadeMux I__8836 (
            .O(N__41049),
            .I(N__41008));
    InMux I__8835 (
            .O(N__41046),
            .I(N__41004));
    InMux I__8834 (
            .O(N__41045),
            .I(N__41001));
    InMux I__8833 (
            .O(N__41044),
            .I(N__40998));
    InMux I__8832 (
            .O(N__41043),
            .I(N__40987));
    InMux I__8831 (
            .O(N__41042),
            .I(N__40987));
    InMux I__8830 (
            .O(N__41041),
            .I(N__40987));
    InMux I__8829 (
            .O(N__41040),
            .I(N__40987));
    InMux I__8828 (
            .O(N__41039),
            .I(N__40987));
    LocalMux I__8827 (
            .O(N__41036),
            .I(N__40984));
    InMux I__8826 (
            .O(N__41035),
            .I(N__40975));
    InMux I__8825 (
            .O(N__41034),
            .I(N__40975));
    InMux I__8824 (
            .O(N__41033),
            .I(N__40975));
    InMux I__8823 (
            .O(N__41032),
            .I(N__40975));
    CascadeMux I__8822 (
            .O(N__41031),
            .I(N__40969));
    CascadeMux I__8821 (
            .O(N__41030),
            .I(N__40966));
    CascadeMux I__8820 (
            .O(N__41029),
            .I(N__40963));
    LocalMux I__8819 (
            .O(N__41026),
            .I(N__40960));
    InMux I__8818 (
            .O(N__41025),
            .I(N__40951));
    InMux I__8817 (
            .O(N__41024),
            .I(N__40951));
    InMux I__8816 (
            .O(N__41023),
            .I(N__40951));
    InMux I__8815 (
            .O(N__41022),
            .I(N__40951));
    LocalMux I__8814 (
            .O(N__41019),
            .I(N__40946));
    LocalMux I__8813 (
            .O(N__41014),
            .I(N__40946));
    InMux I__8812 (
            .O(N__41011),
            .I(N__40943));
    InMux I__8811 (
            .O(N__41008),
            .I(N__40938));
    InMux I__8810 (
            .O(N__41007),
            .I(N__40938));
    LocalMux I__8809 (
            .O(N__41004),
            .I(N__40929));
    LocalMux I__8808 (
            .O(N__41001),
            .I(N__40929));
    LocalMux I__8807 (
            .O(N__40998),
            .I(N__40929));
    LocalMux I__8806 (
            .O(N__40987),
            .I(N__40929));
    Span4Mux_v I__8805 (
            .O(N__40984),
            .I(N__40924));
    LocalMux I__8804 (
            .O(N__40975),
            .I(N__40924));
    InMux I__8803 (
            .O(N__40974),
            .I(N__40917));
    InMux I__8802 (
            .O(N__40973),
            .I(N__40917));
    InMux I__8801 (
            .O(N__40972),
            .I(N__40917));
    InMux I__8800 (
            .O(N__40969),
            .I(N__40910));
    InMux I__8799 (
            .O(N__40966),
            .I(N__40910));
    InMux I__8798 (
            .O(N__40963),
            .I(N__40910));
    Odrv4 I__8797 (
            .O(N__40960),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__8796 (
            .O(N__40951),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__8795 (
            .O(N__40946),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__8794 (
            .O(N__40943),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__8793 (
            .O(N__40938),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__8792 (
            .O(N__40929),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    Odrv4 I__8791 (
            .O(N__40924),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__8790 (
            .O(N__40917),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    LocalMux I__8789 (
            .O(N__40910),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ));
    CascadeMux I__8788 (
            .O(N__40891),
            .I(elapsed_time_ns_1_RNI9865M1_0_17_cascade_));
    InMux I__8787 (
            .O(N__40888),
            .I(N__40885));
    LocalMux I__8786 (
            .O(N__40885),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ));
    InMux I__8785 (
            .O(N__40882),
            .I(N__40879));
    LocalMux I__8784 (
            .O(N__40879),
            .I(N__40876));
    Span4Mux_v I__8783 (
            .O(N__40876),
            .I(N__40873));
    Odrv4 I__8782 (
            .O(N__40873),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ));
    InMux I__8781 (
            .O(N__40870),
            .I(N__40867));
    LocalMux I__8780 (
            .O(N__40867),
            .I(N__40864));
    Odrv4 I__8779 (
            .O(N__40864),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5 ));
    InMux I__8778 (
            .O(N__40861),
            .I(N__40858));
    LocalMux I__8777 (
            .O(N__40858),
            .I(N__40853));
    InMux I__8776 (
            .O(N__40857),
            .I(N__40848));
    InMux I__8775 (
            .O(N__40856),
            .I(N__40848));
    Odrv4 I__8774 (
            .O(N__40853),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lt31_0_2 ));
    LocalMux I__8773 (
            .O(N__40848),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lt31_0_2 ));
    CascadeMux I__8772 (
            .O(N__40843),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4_cascade_ ));
    CascadeMux I__8771 (
            .O(N__40840),
            .I(N__40836));
    InMux I__8770 (
            .O(N__40839),
            .I(N__40832));
    InMux I__8769 (
            .O(N__40836),
            .I(N__40827));
    InMux I__8768 (
            .O(N__40835),
            .I(N__40827));
    LocalMux I__8767 (
            .O(N__40832),
            .I(\delay_measurement_inst.delay_tr_timer.N_358 ));
    LocalMux I__8766 (
            .O(N__40827),
            .I(\delay_measurement_inst.delay_tr_timer.N_358 ));
    InMux I__8765 (
            .O(N__40822),
            .I(N__40810));
    InMux I__8764 (
            .O(N__40821),
            .I(N__40810));
    InMux I__8763 (
            .O(N__40820),
            .I(N__40807));
    InMux I__8762 (
            .O(N__40819),
            .I(N__40804));
    CascadeMux I__8761 (
            .O(N__40818),
            .I(N__40801));
    CascadeMux I__8760 (
            .O(N__40817),
            .I(N__40798));
    CascadeMux I__8759 (
            .O(N__40816),
            .I(N__40795));
    CascadeMux I__8758 (
            .O(N__40815),
            .I(N__40792));
    LocalMux I__8757 (
            .O(N__40810),
            .I(N__40789));
    LocalMux I__8756 (
            .O(N__40807),
            .I(N__40771));
    LocalMux I__8755 (
            .O(N__40804),
            .I(N__40771));
    InMux I__8754 (
            .O(N__40801),
            .I(N__40768));
    InMux I__8753 (
            .O(N__40798),
            .I(N__40761));
    InMux I__8752 (
            .O(N__40795),
            .I(N__40761));
    InMux I__8751 (
            .O(N__40792),
            .I(N__40761));
    Span4Mux_v I__8750 (
            .O(N__40789),
            .I(N__40758));
    InMux I__8749 (
            .O(N__40788),
            .I(N__40755));
    InMux I__8748 (
            .O(N__40787),
            .I(N__40750));
    InMux I__8747 (
            .O(N__40786),
            .I(N__40750));
    InMux I__8746 (
            .O(N__40785),
            .I(N__40745));
    InMux I__8745 (
            .O(N__40784),
            .I(N__40745));
    InMux I__8744 (
            .O(N__40783),
            .I(N__40740));
    InMux I__8743 (
            .O(N__40782),
            .I(N__40740));
    InMux I__8742 (
            .O(N__40781),
            .I(N__40733));
    InMux I__8741 (
            .O(N__40780),
            .I(N__40733));
    InMux I__8740 (
            .O(N__40779),
            .I(N__40733));
    InMux I__8739 (
            .O(N__40778),
            .I(N__40726));
    InMux I__8738 (
            .O(N__40777),
            .I(N__40726));
    InMux I__8737 (
            .O(N__40776),
            .I(N__40726));
    Odrv4 I__8736 (
            .O(N__40771),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8735 (
            .O(N__40768),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8734 (
            .O(N__40761),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    Odrv4 I__8733 (
            .O(N__40758),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8732 (
            .O(N__40755),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8731 (
            .O(N__40750),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8730 (
            .O(N__40745),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8729 (
            .O(N__40740),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8728 (
            .O(N__40733),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    LocalMux I__8727 (
            .O(N__40726),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ));
    InMux I__8726 (
            .O(N__40705),
            .I(N__40702));
    LocalMux I__8725 (
            .O(N__40702),
            .I(\delay_measurement_inst.delay_tr_timer.N_354 ));
    CascadeMux I__8724 (
            .O(N__40699),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ));
    InMux I__8723 (
            .O(N__40696),
            .I(N__40693));
    LocalMux I__8722 (
            .O(N__40693),
            .I(N__40689));
    InMux I__8721 (
            .O(N__40692),
            .I(N__40686));
    Span4Mux_v I__8720 (
            .O(N__40689),
            .I(N__40681));
    LocalMux I__8719 (
            .O(N__40686),
            .I(N__40678));
    InMux I__8718 (
            .O(N__40685),
            .I(N__40675));
    InMux I__8717 (
            .O(N__40684),
            .I(N__40671));
    Span4Mux_h I__8716 (
            .O(N__40681),
            .I(N__40668));
    Span4Mux_v I__8715 (
            .O(N__40678),
            .I(N__40663));
    LocalMux I__8714 (
            .O(N__40675),
            .I(N__40663));
    InMux I__8713 (
            .O(N__40674),
            .I(N__40660));
    LocalMux I__8712 (
            .O(N__40671),
            .I(elapsed_time_ns_1_RNIK8NQL1_0_3));
    Odrv4 I__8711 (
            .O(N__40668),
            .I(elapsed_time_ns_1_RNIK8NQL1_0_3));
    Odrv4 I__8710 (
            .O(N__40663),
            .I(elapsed_time_ns_1_RNIK8NQL1_0_3));
    LocalMux I__8709 (
            .O(N__40660),
            .I(elapsed_time_ns_1_RNIK8NQL1_0_3));
    InMux I__8708 (
            .O(N__40651),
            .I(N__40648));
    LocalMux I__8707 (
            .O(N__40648),
            .I(N__40645));
    Odrv4 I__8706 (
            .O(N__40645),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6 ));
    CascadeMux I__8705 (
            .O(N__40642),
            .I(N__40639));
    InMux I__8704 (
            .O(N__40639),
            .I(N__40635));
    InMux I__8703 (
            .O(N__40638),
            .I(N__40631));
    LocalMux I__8702 (
            .O(N__40635),
            .I(N__40627));
    InMux I__8701 (
            .O(N__40634),
            .I(N__40624));
    LocalMux I__8700 (
            .O(N__40631),
            .I(N__40621));
    InMux I__8699 (
            .O(N__40630),
            .I(N__40618));
    Span4Mux_v I__8698 (
            .O(N__40627),
            .I(N__40613));
    LocalMux I__8697 (
            .O(N__40624),
            .I(N__40613));
    Odrv4 I__8696 (
            .O(N__40621),
            .I(elapsed_time_ns_1_RNINBNQL1_0_6));
    LocalMux I__8695 (
            .O(N__40618),
            .I(elapsed_time_ns_1_RNINBNQL1_0_6));
    Odrv4 I__8694 (
            .O(N__40613),
            .I(elapsed_time_ns_1_RNINBNQL1_0_6));
    InMux I__8693 (
            .O(N__40606),
            .I(N__40603));
    LocalMux I__8692 (
            .O(N__40603),
            .I(\delay_measurement_inst.delay_tr_timer.N_353 ));
    CascadeMux I__8691 (
            .O(N__40600),
            .I(elapsed_time_ns_1_RNITCIF91_0_23_cascade_));
    CascadeMux I__8690 (
            .O(N__40597),
            .I(N__40594));
    InMux I__8689 (
            .O(N__40594),
            .I(N__40591));
    LocalMux I__8688 (
            .O(N__40591),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ));
    CascadeMux I__8687 (
            .O(N__40588),
            .I(N__40585));
    InMux I__8686 (
            .O(N__40585),
            .I(N__40581));
    InMux I__8685 (
            .O(N__40584),
            .I(N__40578));
    LocalMux I__8684 (
            .O(N__40581),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    LocalMux I__8683 (
            .O(N__40578),
            .I(elapsed_time_ns_1_RNIUDIF91_0_24));
    CascadeMux I__8682 (
            .O(N__40573),
            .I(\delay_measurement_inst.delay_tr_timer.N_379_cascade_ ));
    CascadeMux I__8681 (
            .O(N__40570),
            .I(\delay_measurement_inst.delay_tr9_cascade_ ));
    CascadeMux I__8680 (
            .O(N__40567),
            .I(N__40564));
    InMux I__8679 (
            .O(N__40564),
            .I(N__40560));
    InMux I__8678 (
            .O(N__40563),
            .I(N__40557));
    LocalMux I__8677 (
            .O(N__40560),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    LocalMux I__8676 (
            .O(N__40557),
            .I(elapsed_time_ns_1_RNIRBJF91_0_30));
    InMux I__8675 (
            .O(N__40552),
            .I(N__40545));
    InMux I__8674 (
            .O(N__40551),
            .I(N__40545));
    InMux I__8673 (
            .O(N__40550),
            .I(N__40542));
    LocalMux I__8672 (
            .O(N__40545),
            .I(N__40539));
    LocalMux I__8671 (
            .O(N__40542),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv12 I__8670 (
            .O(N__40539),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__8669 (
            .O(N__40534),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__8668 (
            .O(N__40531),
            .I(N__40527));
    CascadeMux I__8667 (
            .O(N__40530),
            .I(N__40524));
    InMux I__8666 (
            .O(N__40527),
            .I(N__40518));
    InMux I__8665 (
            .O(N__40524),
            .I(N__40518));
    InMux I__8664 (
            .O(N__40523),
            .I(N__40515));
    LocalMux I__8663 (
            .O(N__40518),
            .I(N__40512));
    LocalMux I__8662 (
            .O(N__40515),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv12 I__8661 (
            .O(N__40512),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__8660 (
            .O(N__40507),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    CascadeMux I__8659 (
            .O(N__40504),
            .I(N__40501));
    InMux I__8658 (
            .O(N__40501),
            .I(N__40497));
    InMux I__8657 (
            .O(N__40500),
            .I(N__40494));
    LocalMux I__8656 (
            .O(N__40497),
            .I(N__40491));
    LocalMux I__8655 (
            .O(N__40494),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv12 I__8654 (
            .O(N__40491),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__8653 (
            .O(N__40486),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__8652 (
            .O(N__40483),
            .I(N__40467));
    InMux I__8651 (
            .O(N__40482),
            .I(N__40467));
    InMux I__8650 (
            .O(N__40481),
            .I(N__40467));
    InMux I__8649 (
            .O(N__40480),
            .I(N__40467));
    InMux I__8648 (
            .O(N__40479),
            .I(N__40444));
    InMux I__8647 (
            .O(N__40478),
            .I(N__40444));
    InMux I__8646 (
            .O(N__40477),
            .I(N__40444));
    InMux I__8645 (
            .O(N__40476),
            .I(N__40444));
    LocalMux I__8644 (
            .O(N__40467),
            .I(N__40437));
    InMux I__8643 (
            .O(N__40466),
            .I(N__40432));
    InMux I__8642 (
            .O(N__40465),
            .I(N__40432));
    InMux I__8641 (
            .O(N__40464),
            .I(N__40423));
    InMux I__8640 (
            .O(N__40463),
            .I(N__40423));
    InMux I__8639 (
            .O(N__40462),
            .I(N__40423));
    InMux I__8638 (
            .O(N__40461),
            .I(N__40423));
    InMux I__8637 (
            .O(N__40460),
            .I(N__40414));
    InMux I__8636 (
            .O(N__40459),
            .I(N__40414));
    InMux I__8635 (
            .O(N__40458),
            .I(N__40414));
    InMux I__8634 (
            .O(N__40457),
            .I(N__40414));
    InMux I__8633 (
            .O(N__40456),
            .I(N__40405));
    InMux I__8632 (
            .O(N__40455),
            .I(N__40405));
    InMux I__8631 (
            .O(N__40454),
            .I(N__40405));
    InMux I__8630 (
            .O(N__40453),
            .I(N__40405));
    LocalMux I__8629 (
            .O(N__40444),
            .I(N__40398));
    InMux I__8628 (
            .O(N__40443),
            .I(N__40389));
    InMux I__8627 (
            .O(N__40442),
            .I(N__40389));
    InMux I__8626 (
            .O(N__40441),
            .I(N__40389));
    InMux I__8625 (
            .O(N__40440),
            .I(N__40389));
    Span4Mux_v I__8624 (
            .O(N__40437),
            .I(N__40382));
    LocalMux I__8623 (
            .O(N__40432),
            .I(N__40382));
    LocalMux I__8622 (
            .O(N__40423),
            .I(N__40382));
    LocalMux I__8621 (
            .O(N__40414),
            .I(N__40379));
    LocalMux I__8620 (
            .O(N__40405),
            .I(N__40376));
    InMux I__8619 (
            .O(N__40404),
            .I(N__40367));
    InMux I__8618 (
            .O(N__40403),
            .I(N__40367));
    InMux I__8617 (
            .O(N__40402),
            .I(N__40367));
    InMux I__8616 (
            .O(N__40401),
            .I(N__40367));
    Span4Mux_v I__8615 (
            .O(N__40398),
            .I(N__40358));
    LocalMux I__8614 (
            .O(N__40389),
            .I(N__40358));
    Span4Mux_v I__8613 (
            .O(N__40382),
            .I(N__40358));
    Span4Mux_v I__8612 (
            .O(N__40379),
            .I(N__40358));
    Span4Mux_v I__8611 (
            .O(N__40376),
            .I(N__40353));
    LocalMux I__8610 (
            .O(N__40367),
            .I(N__40353));
    Span4Mux_h I__8609 (
            .O(N__40358),
            .I(N__40348));
    Span4Mux_h I__8608 (
            .O(N__40353),
            .I(N__40348));
    Odrv4 I__8607 (
            .O(N__40348),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__8606 (
            .O(N__40345),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__8605 (
            .O(N__40342),
            .I(N__40338));
    InMux I__8604 (
            .O(N__40341),
            .I(N__40335));
    LocalMux I__8603 (
            .O(N__40338),
            .I(N__40332));
    LocalMux I__8602 (
            .O(N__40335),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv12 I__8601 (
            .O(N__40332),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CEMux I__8600 (
            .O(N__40327),
            .I(N__40322));
    CEMux I__8599 (
            .O(N__40326),
            .I(N__40319));
    CEMux I__8598 (
            .O(N__40325),
            .I(N__40315));
    LocalMux I__8597 (
            .O(N__40322),
            .I(N__40310));
    LocalMux I__8596 (
            .O(N__40319),
            .I(N__40310));
    CEMux I__8595 (
            .O(N__40318),
            .I(N__40307));
    LocalMux I__8594 (
            .O(N__40315),
            .I(N__40304));
    Span4Mux_v I__8593 (
            .O(N__40310),
            .I(N__40301));
    LocalMux I__8592 (
            .O(N__40307),
            .I(N__40298));
    Span4Mux_v I__8591 (
            .O(N__40304),
            .I(N__40291));
    Span4Mux_h I__8590 (
            .O(N__40301),
            .I(N__40291));
    Span4Mux_h I__8589 (
            .O(N__40298),
            .I(N__40291));
    Span4Mux_h I__8588 (
            .O(N__40291),
            .I(N__40288));
    Odrv4 I__8587 (
            .O(N__40288),
            .I(\delay_measurement_inst.delay_hc_timer.N_398_i ));
    InMux I__8586 (
            .O(N__40285),
            .I(N__40282));
    LocalMux I__8585 (
            .O(N__40282),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20));
    InMux I__8584 (
            .O(N__40279),
            .I(N__40275));
    InMux I__8583 (
            .O(N__40278),
            .I(N__40272));
    LocalMux I__8582 (
            .O(N__40275),
            .I(elapsed_time_ns_1_RNIRAIF91_0_21));
    LocalMux I__8581 (
            .O(N__40272),
            .I(elapsed_time_ns_1_RNIRAIF91_0_21));
    CascadeMux I__8580 (
            .O(N__40267),
            .I(elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_));
    InMux I__8579 (
            .O(N__40264),
            .I(N__40258));
    InMux I__8578 (
            .O(N__40263),
            .I(N__40258));
    LocalMux I__8577 (
            .O(N__40258),
            .I(elapsed_time_ns_1_RNI3JIF91_0_29));
    InMux I__8576 (
            .O(N__40255),
            .I(N__40252));
    LocalMux I__8575 (
            .O(N__40252),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15 ));
    InMux I__8574 (
            .O(N__40249),
            .I(N__40246));
    LocalMux I__8573 (
            .O(N__40246),
            .I(elapsed_time_ns_1_RNITCIF91_0_23));
    InMux I__8572 (
            .O(N__40243),
            .I(N__40240));
    LocalMux I__8571 (
            .O(N__40240),
            .I(N__40235));
    InMux I__8570 (
            .O(N__40239),
            .I(N__40232));
    InMux I__8569 (
            .O(N__40238),
            .I(N__40229));
    Span4Mux_h I__8568 (
            .O(N__40235),
            .I(N__40226));
    LocalMux I__8567 (
            .O(N__40232),
            .I(N__40223));
    LocalMux I__8566 (
            .O(N__40229),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__8565 (
            .O(N__40226),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv12 I__8564 (
            .O(N__40223),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__8563 (
            .O(N__40216),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    CascadeMux I__8562 (
            .O(N__40213),
            .I(N__40210));
    InMux I__8561 (
            .O(N__40210),
            .I(N__40206));
    InMux I__8560 (
            .O(N__40209),
            .I(N__40203));
    LocalMux I__8559 (
            .O(N__40206),
            .I(N__40197));
    LocalMux I__8558 (
            .O(N__40203),
            .I(N__40197));
    InMux I__8557 (
            .O(N__40202),
            .I(N__40194));
    Span4Mux_h I__8556 (
            .O(N__40197),
            .I(N__40191));
    LocalMux I__8555 (
            .O(N__40194),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__8554 (
            .O(N__40191),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__8553 (
            .O(N__40186),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    CascadeMux I__8552 (
            .O(N__40183),
            .I(N__40179));
    CascadeMux I__8551 (
            .O(N__40182),
            .I(N__40176));
    InMux I__8550 (
            .O(N__40179),
            .I(N__40170));
    InMux I__8549 (
            .O(N__40176),
            .I(N__40170));
    InMux I__8548 (
            .O(N__40175),
            .I(N__40167));
    LocalMux I__8547 (
            .O(N__40170),
            .I(N__40164));
    LocalMux I__8546 (
            .O(N__40167),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv12 I__8545 (
            .O(N__40164),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__8544 (
            .O(N__40159),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__8543 (
            .O(N__40156),
            .I(N__40149));
    InMux I__8542 (
            .O(N__40155),
            .I(N__40149));
    InMux I__8541 (
            .O(N__40154),
            .I(N__40146));
    LocalMux I__8540 (
            .O(N__40149),
            .I(N__40143));
    LocalMux I__8539 (
            .O(N__40146),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv12 I__8538 (
            .O(N__40143),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__8537 (
            .O(N__40138),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__8536 (
            .O(N__40135),
            .I(N__40132));
    InMux I__8535 (
            .O(N__40132),
            .I(N__40127));
    InMux I__8534 (
            .O(N__40131),
            .I(N__40124));
    InMux I__8533 (
            .O(N__40130),
            .I(N__40121));
    LocalMux I__8532 (
            .O(N__40127),
            .I(N__40116));
    LocalMux I__8531 (
            .O(N__40124),
            .I(N__40116));
    LocalMux I__8530 (
            .O(N__40121),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv12 I__8529 (
            .O(N__40116),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__8528 (
            .O(N__40111),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    CascadeMux I__8527 (
            .O(N__40108),
            .I(N__40104));
    CascadeMux I__8526 (
            .O(N__40107),
            .I(N__40101));
    InMux I__8525 (
            .O(N__40104),
            .I(N__40096));
    InMux I__8524 (
            .O(N__40101),
            .I(N__40096));
    LocalMux I__8523 (
            .O(N__40096),
            .I(N__40092));
    InMux I__8522 (
            .O(N__40095),
            .I(N__40089));
    Span4Mux_v I__8521 (
            .O(N__40092),
            .I(N__40086));
    LocalMux I__8520 (
            .O(N__40089),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__8519 (
            .O(N__40086),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__8518 (
            .O(N__40081),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__8517 (
            .O(N__40078),
            .I(N__40071));
    InMux I__8516 (
            .O(N__40077),
            .I(N__40071));
    InMux I__8515 (
            .O(N__40076),
            .I(N__40068));
    LocalMux I__8514 (
            .O(N__40071),
            .I(N__40065));
    LocalMux I__8513 (
            .O(N__40068),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv12 I__8512 (
            .O(N__40065),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__8511 (
            .O(N__40060),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__8510 (
            .O(N__40057),
            .I(N__40054));
    InMux I__8509 (
            .O(N__40054),
            .I(N__40051));
    LocalMux I__8508 (
            .O(N__40051),
            .I(N__40046));
    InMux I__8507 (
            .O(N__40050),
            .I(N__40043));
    InMux I__8506 (
            .O(N__40049),
            .I(N__40040));
    Span4Mux_h I__8505 (
            .O(N__40046),
            .I(N__40037));
    LocalMux I__8504 (
            .O(N__40043),
            .I(N__40034));
    LocalMux I__8503 (
            .O(N__40040),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__8502 (
            .O(N__40037),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv12 I__8501 (
            .O(N__40034),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__8500 (
            .O(N__40027),
            .I(bfn_15_24_0_));
    InMux I__8499 (
            .O(N__40024),
            .I(N__40020));
    CascadeMux I__8498 (
            .O(N__40023),
            .I(N__40017));
    LocalMux I__8497 (
            .O(N__40020),
            .I(N__40013));
    InMux I__8496 (
            .O(N__40017),
            .I(N__40010));
    InMux I__8495 (
            .O(N__40016),
            .I(N__40007));
    Span4Mux_h I__8494 (
            .O(N__40013),
            .I(N__40004));
    LocalMux I__8493 (
            .O(N__40010),
            .I(N__40001));
    LocalMux I__8492 (
            .O(N__40007),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__8491 (
            .O(N__40004),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv12 I__8490 (
            .O(N__40001),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__8489 (
            .O(N__39994),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__8488 (
            .O(N__39991),
            .I(N__39988));
    InMux I__8487 (
            .O(N__39988),
            .I(N__39984));
    InMux I__8486 (
            .O(N__39987),
            .I(N__39981));
    LocalMux I__8485 (
            .O(N__39984),
            .I(N__39975));
    LocalMux I__8484 (
            .O(N__39981),
            .I(N__39975));
    InMux I__8483 (
            .O(N__39980),
            .I(N__39972));
    Span4Mux_v I__8482 (
            .O(N__39975),
            .I(N__39969));
    LocalMux I__8481 (
            .O(N__39972),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__8480 (
            .O(N__39969),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__8479 (
            .O(N__39964),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__8478 (
            .O(N__39961),
            .I(N__39955));
    InMux I__8477 (
            .O(N__39960),
            .I(N__39955));
    LocalMux I__8476 (
            .O(N__39955),
            .I(N__39951));
    InMux I__8475 (
            .O(N__39954),
            .I(N__39948));
    Span4Mux_h I__8474 (
            .O(N__39951),
            .I(N__39945));
    LocalMux I__8473 (
            .O(N__39948),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__8472 (
            .O(N__39945),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__8471 (
            .O(N__39940),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__8470 (
            .O(N__39937),
            .I(N__39931));
    InMux I__8469 (
            .O(N__39936),
            .I(N__39931));
    LocalMux I__8468 (
            .O(N__39931),
            .I(N__39927));
    InMux I__8467 (
            .O(N__39930),
            .I(N__39924));
    Span4Mux_h I__8466 (
            .O(N__39927),
            .I(N__39921));
    LocalMux I__8465 (
            .O(N__39924),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__8464 (
            .O(N__39921),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__8463 (
            .O(N__39916),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    CascadeMux I__8462 (
            .O(N__39913),
            .I(N__39909));
    CascadeMux I__8461 (
            .O(N__39912),
            .I(N__39906));
    InMux I__8460 (
            .O(N__39909),
            .I(N__39901));
    InMux I__8459 (
            .O(N__39906),
            .I(N__39901));
    LocalMux I__8458 (
            .O(N__39901),
            .I(N__39897));
    InMux I__8457 (
            .O(N__39900),
            .I(N__39894));
    Span4Mux_v I__8456 (
            .O(N__39897),
            .I(N__39891));
    LocalMux I__8455 (
            .O(N__39894),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__8454 (
            .O(N__39891),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__8453 (
            .O(N__39886),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    CascadeMux I__8452 (
            .O(N__39883),
            .I(N__39879));
    CascadeMux I__8451 (
            .O(N__39882),
            .I(N__39876));
    InMux I__8450 (
            .O(N__39879),
            .I(N__39871));
    InMux I__8449 (
            .O(N__39876),
            .I(N__39871));
    LocalMux I__8448 (
            .O(N__39871),
            .I(N__39867));
    InMux I__8447 (
            .O(N__39870),
            .I(N__39864));
    Span4Mux_h I__8446 (
            .O(N__39867),
            .I(N__39861));
    LocalMux I__8445 (
            .O(N__39864),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__8444 (
            .O(N__39861),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__8443 (
            .O(N__39856),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    CascadeMux I__8442 (
            .O(N__39853),
            .I(N__39850));
    InMux I__8441 (
            .O(N__39850),
            .I(N__39846));
    InMux I__8440 (
            .O(N__39849),
            .I(N__39843));
    LocalMux I__8439 (
            .O(N__39846),
            .I(N__39837));
    LocalMux I__8438 (
            .O(N__39843),
            .I(N__39837));
    InMux I__8437 (
            .O(N__39842),
            .I(N__39834));
    Span4Mux_v I__8436 (
            .O(N__39837),
            .I(N__39831));
    LocalMux I__8435 (
            .O(N__39834),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__8434 (
            .O(N__39831),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__8433 (
            .O(N__39826),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    CascadeMux I__8432 (
            .O(N__39823),
            .I(N__39820));
    InMux I__8431 (
            .O(N__39820),
            .I(N__39816));
    InMux I__8430 (
            .O(N__39819),
            .I(N__39813));
    LocalMux I__8429 (
            .O(N__39816),
            .I(N__39807));
    LocalMux I__8428 (
            .O(N__39813),
            .I(N__39807));
    InMux I__8427 (
            .O(N__39812),
            .I(N__39804));
    Span4Mux_v I__8426 (
            .O(N__39807),
            .I(N__39801));
    LocalMux I__8425 (
            .O(N__39804),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__8424 (
            .O(N__39801),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__8423 (
            .O(N__39796),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__8422 (
            .O(N__39793),
            .I(N__39790));
    InMux I__8421 (
            .O(N__39790),
            .I(N__39786));
    InMux I__8420 (
            .O(N__39789),
            .I(N__39783));
    LocalMux I__8419 (
            .O(N__39786),
            .I(N__39779));
    LocalMux I__8418 (
            .O(N__39783),
            .I(N__39776));
    InMux I__8417 (
            .O(N__39782),
            .I(N__39773));
    Span4Mux_v I__8416 (
            .O(N__39779),
            .I(N__39768));
    Span4Mux_v I__8415 (
            .O(N__39776),
            .I(N__39768));
    LocalMux I__8414 (
            .O(N__39773),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__8413 (
            .O(N__39768),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__8412 (
            .O(N__39763),
            .I(bfn_15_23_0_));
    CascadeMux I__8411 (
            .O(N__39760),
            .I(N__39756));
    InMux I__8410 (
            .O(N__39759),
            .I(N__39753));
    InMux I__8409 (
            .O(N__39756),
            .I(N__39750));
    LocalMux I__8408 (
            .O(N__39753),
            .I(N__39747));
    LocalMux I__8407 (
            .O(N__39750),
            .I(N__39743));
    Span4Mux_h I__8406 (
            .O(N__39747),
            .I(N__39740));
    InMux I__8405 (
            .O(N__39746),
            .I(N__39737));
    Span4Mux_h I__8404 (
            .O(N__39743),
            .I(N__39734));
    Odrv4 I__8403 (
            .O(N__39740),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__8402 (
            .O(N__39737),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__8401 (
            .O(N__39734),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__8400 (
            .O(N__39727),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__8399 (
            .O(N__39724),
            .I(N__39717));
    InMux I__8398 (
            .O(N__39723),
            .I(N__39717));
    InMux I__8397 (
            .O(N__39722),
            .I(N__39714));
    LocalMux I__8396 (
            .O(N__39717),
            .I(N__39711));
    LocalMux I__8395 (
            .O(N__39714),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv12 I__8394 (
            .O(N__39711),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__8393 (
            .O(N__39706),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__8392 (
            .O(N__39703),
            .I(N__39697));
    InMux I__8391 (
            .O(N__39702),
            .I(N__39697));
    LocalMux I__8390 (
            .O(N__39697),
            .I(N__39693));
    InMux I__8389 (
            .O(N__39696),
            .I(N__39690));
    Span4Mux_v I__8388 (
            .O(N__39693),
            .I(N__39687));
    LocalMux I__8387 (
            .O(N__39690),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__8386 (
            .O(N__39687),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__8385 (
            .O(N__39682),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__8384 (
            .O(N__39679),
            .I(N__39675));
    InMux I__8383 (
            .O(N__39678),
            .I(N__39671));
    InMux I__8382 (
            .O(N__39675),
            .I(N__39668));
    InMux I__8381 (
            .O(N__39674),
            .I(N__39665));
    LocalMux I__8380 (
            .O(N__39671),
            .I(N__39660));
    LocalMux I__8379 (
            .O(N__39668),
            .I(N__39660));
    LocalMux I__8378 (
            .O(N__39665),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv12 I__8377 (
            .O(N__39660),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__8376 (
            .O(N__39655),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__8375 (
            .O(N__39652),
            .I(N__39648));
    CascadeMux I__8374 (
            .O(N__39651),
            .I(N__39645));
    InMux I__8373 (
            .O(N__39648),
            .I(N__39640));
    InMux I__8372 (
            .O(N__39645),
            .I(N__39640));
    LocalMux I__8371 (
            .O(N__39640),
            .I(N__39636));
    InMux I__8370 (
            .O(N__39639),
            .I(N__39633));
    Span4Mux_h I__8369 (
            .O(N__39636),
            .I(N__39630));
    LocalMux I__8368 (
            .O(N__39633),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__8367 (
            .O(N__39630),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__8366 (
            .O(N__39625),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    CascadeMux I__8365 (
            .O(N__39622),
            .I(N__39618));
    CascadeMux I__8364 (
            .O(N__39621),
            .I(N__39615));
    InMux I__8363 (
            .O(N__39618),
            .I(N__39610));
    InMux I__8362 (
            .O(N__39615),
            .I(N__39610));
    LocalMux I__8361 (
            .O(N__39610),
            .I(N__39606));
    InMux I__8360 (
            .O(N__39609),
            .I(N__39603));
    Span4Mux_v I__8359 (
            .O(N__39606),
            .I(N__39600));
    LocalMux I__8358 (
            .O(N__39603),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__8357 (
            .O(N__39600),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__8356 (
            .O(N__39595),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    CascadeMux I__8355 (
            .O(N__39592),
            .I(N__39589));
    InMux I__8354 (
            .O(N__39589),
            .I(N__39585));
    InMux I__8353 (
            .O(N__39588),
            .I(N__39582));
    LocalMux I__8352 (
            .O(N__39585),
            .I(N__39576));
    LocalMux I__8351 (
            .O(N__39582),
            .I(N__39576));
    InMux I__8350 (
            .O(N__39581),
            .I(N__39573));
    Span4Mux_v I__8349 (
            .O(N__39576),
            .I(N__39570));
    LocalMux I__8348 (
            .O(N__39573),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__8347 (
            .O(N__39570),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__8346 (
            .O(N__39565),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    CascadeMux I__8345 (
            .O(N__39562),
            .I(N__39559));
    InMux I__8344 (
            .O(N__39559),
            .I(N__39556));
    LocalMux I__8343 (
            .O(N__39556),
            .I(N__39551));
    InMux I__8342 (
            .O(N__39555),
            .I(N__39548));
    InMux I__8341 (
            .O(N__39554),
            .I(N__39545));
    Span4Mux_h I__8340 (
            .O(N__39551),
            .I(N__39542));
    LocalMux I__8339 (
            .O(N__39548),
            .I(N__39539));
    LocalMux I__8338 (
            .O(N__39545),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__8337 (
            .O(N__39542),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv12 I__8336 (
            .O(N__39539),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__8335 (
            .O(N__39532),
            .I(bfn_15_22_0_));
    InMux I__8334 (
            .O(N__39529),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__8333 (
            .O(N__39526),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__8332 (
            .O(N__39523),
            .I(bfn_15_20_0_));
    InMux I__8331 (
            .O(N__39520),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__8330 (
            .O(N__39517),
            .I(N__39513));
    InMux I__8329 (
            .O(N__39516),
            .I(N__39510));
    LocalMux I__8328 (
            .O(N__39513),
            .I(N__39507));
    LocalMux I__8327 (
            .O(N__39510),
            .I(N__39504));
    Span4Mux_v I__8326 (
            .O(N__39507),
            .I(N__39499));
    Span4Mux_h I__8325 (
            .O(N__39504),
            .I(N__39499));
    Odrv4 I__8324 (
            .O(N__39499),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__8323 (
            .O(N__39496),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    CascadeMux I__8322 (
            .O(N__39493),
            .I(N__39490));
    InMux I__8321 (
            .O(N__39490),
            .I(N__39486));
    InMux I__8320 (
            .O(N__39489),
            .I(N__39483));
    LocalMux I__8319 (
            .O(N__39486),
            .I(N__39480));
    LocalMux I__8318 (
            .O(N__39483),
            .I(N__39477));
    Span4Mux_h I__8317 (
            .O(N__39480),
            .I(N__39474));
    Odrv12 I__8316 (
            .O(N__39477),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__8315 (
            .O(N__39474),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__8314 (
            .O(N__39469),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__8313 (
            .O(N__39466),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__8312 (
            .O(N__39463),
            .I(N__39460));
    LocalMux I__8311 (
            .O(N__39460),
            .I(N__39457));
    Span4Mux_h I__8310 (
            .O(N__39457),
            .I(N__39454));
    Odrv4 I__8309 (
            .O(N__39454),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    CEMux I__8308 (
            .O(N__39451),
            .I(N__39436));
    CEMux I__8307 (
            .O(N__39450),
            .I(N__39436));
    CEMux I__8306 (
            .O(N__39449),
            .I(N__39436));
    CEMux I__8305 (
            .O(N__39448),
            .I(N__39436));
    CEMux I__8304 (
            .O(N__39447),
            .I(N__39436));
    GlobalMux I__8303 (
            .O(N__39436),
            .I(N__39433));
    gio2CtrlBuf I__8302 (
            .O(N__39433),
            .I(\delay_measurement_inst.delay_hc_timer.N_397_i_g ));
    CascadeMux I__8301 (
            .O(N__39430),
            .I(N__39427));
    InMux I__8300 (
            .O(N__39427),
            .I(N__39424));
    LocalMux I__8299 (
            .O(N__39424),
            .I(N__39419));
    InMux I__8298 (
            .O(N__39423),
            .I(N__39416));
    InMux I__8297 (
            .O(N__39422),
            .I(N__39413));
    Span4Mux_h I__8296 (
            .O(N__39419),
            .I(N__39410));
    LocalMux I__8295 (
            .O(N__39416),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__8294 (
            .O(N__39413),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv4 I__8293 (
            .O(N__39410),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__8292 (
            .O(N__39403),
            .I(bfn_15_21_0_));
    InMux I__8291 (
            .O(N__39400),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__8290 (
            .O(N__39397),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__8289 (
            .O(N__39394),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__8288 (
            .O(N__39391),
            .I(bfn_15_19_0_));
    InMux I__8287 (
            .O(N__39388),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__8286 (
            .O(N__39385),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__8285 (
            .O(N__39382),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__8284 (
            .O(N__39379),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__8283 (
            .O(N__39376),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__8282 (
            .O(N__39373),
            .I(N__39367));
    InMux I__8281 (
            .O(N__39372),
            .I(N__39367));
    LocalMux I__8280 (
            .O(N__39367),
            .I(N__39364));
    Odrv4 I__8279 (
            .O(N__39364),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__8278 (
            .O(N__39361),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__8277 (
            .O(N__39358),
            .I(N__39352));
    InMux I__8276 (
            .O(N__39357),
            .I(N__39352));
    LocalMux I__8275 (
            .O(N__39352),
            .I(N__39349));
    Odrv12 I__8274 (
            .O(N__39349),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__8273 (
            .O(N__39346),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__8272 (
            .O(N__39343),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__8271 (
            .O(N__39340),
            .I(N__39336));
    InMux I__8270 (
            .O(N__39339),
            .I(N__39333));
    LocalMux I__8269 (
            .O(N__39336),
            .I(N__39330));
    LocalMux I__8268 (
            .O(N__39333),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    Odrv4 I__8267 (
            .O(N__39330),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__8266 (
            .O(N__39325),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__8265 (
            .O(N__39322),
            .I(bfn_15_18_0_));
    InMux I__8264 (
            .O(N__39319),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__8263 (
            .O(N__39316),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__8262 (
            .O(N__39313),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__8261 (
            .O(N__39310),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__8260 (
            .O(N__39307),
            .I(N__39304));
    LocalMux I__8259 (
            .O(N__39304),
            .I(N__39300));
    InMux I__8258 (
            .O(N__39303),
            .I(N__39297));
    Span4Mux_h I__8257 (
            .O(N__39300),
            .I(N__39293));
    LocalMux I__8256 (
            .O(N__39297),
            .I(N__39290));
    CascadeMux I__8255 (
            .O(N__39296),
            .I(N__39287));
    Span4Mux_h I__8254 (
            .O(N__39293),
            .I(N__39284));
    Span4Mux_v I__8253 (
            .O(N__39290),
            .I(N__39281));
    InMux I__8252 (
            .O(N__39287),
            .I(N__39278));
    Odrv4 I__8251 (
            .O(N__39284),
            .I(elapsed_time_ns_1_RNILGKEE1_0_4));
    Odrv4 I__8250 (
            .O(N__39281),
            .I(elapsed_time_ns_1_RNILGKEE1_0_4));
    LocalMux I__8249 (
            .O(N__39278),
            .I(elapsed_time_ns_1_RNILGKEE1_0_4));
    CascadeMux I__8248 (
            .O(N__39271),
            .I(elapsed_time_ns_1_RNILGKEE1_0_4_cascade_));
    InMux I__8247 (
            .O(N__39268),
            .I(N__39265));
    LocalMux I__8246 (
            .O(N__39265),
            .I(N__39262));
    Odrv4 I__8245 (
            .O(N__39262),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2 ));
    InMux I__8244 (
            .O(N__39259),
            .I(N__39253));
    InMux I__8243 (
            .O(N__39258),
            .I(N__39253));
    LocalMux I__8242 (
            .O(N__39253),
            .I(elapsed_time_ns_1_RNI4GU8E1_0_21));
    InMux I__8241 (
            .O(N__39250),
            .I(N__39244));
    InMux I__8240 (
            .O(N__39249),
            .I(N__39244));
    LocalMux I__8239 (
            .O(N__39244),
            .I(elapsed_time_ns_1_RNICOU8E1_0_29));
    InMux I__8238 (
            .O(N__39241),
            .I(N__39237));
    InMux I__8237 (
            .O(N__39240),
            .I(N__39234));
    LocalMux I__8236 (
            .O(N__39237),
            .I(N__39229));
    LocalMux I__8235 (
            .O(N__39234),
            .I(N__39229));
    Span4Mux_h I__8234 (
            .O(N__39229),
            .I(N__39226));
    Odrv4 I__8233 (
            .O(N__39226),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__8232 (
            .O(N__39223),
            .I(N__39220));
    LocalMux I__8231 (
            .O(N__39220),
            .I(N__39216));
    InMux I__8230 (
            .O(N__39219),
            .I(N__39213));
    Span4Mux_h I__8229 (
            .O(N__39216),
            .I(N__39210));
    LocalMux I__8228 (
            .O(N__39213),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__8227 (
            .O(N__39210),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__8226 (
            .O(N__39205),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__8225 (
            .O(N__39202),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__8224 (
            .O(N__39199),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__8223 (
            .O(N__39196),
            .I(N__39193));
    LocalMux I__8222 (
            .O(N__39193),
            .I(N__39190));
    Span4Mux_h I__8221 (
            .O(N__39190),
            .I(N__39187));
    Odrv4 I__8220 (
            .O(N__39187),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df22 ));
    InMux I__8219 (
            .O(N__39184),
            .I(N__39181));
    LocalMux I__8218 (
            .O(N__39181),
            .I(N__39178));
    Span4Mux_v I__8217 (
            .O(N__39178),
            .I(N__39175));
    Odrv4 I__8216 (
            .O(N__39175),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df24 ));
    InMux I__8215 (
            .O(N__39172),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ));
    InMux I__8214 (
            .O(N__39169),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    CascadeMux I__8213 (
            .O(N__39166),
            .I(N__39162));
    InMux I__8212 (
            .O(N__39165),
            .I(N__39157));
    InMux I__8211 (
            .O(N__39162),
            .I(N__39157));
    LocalMux I__8210 (
            .O(N__39157),
            .I(elapsed_time_ns_1_RNI4HV8E1_0_30));
    CascadeMux I__8209 (
            .O(N__39154),
            .I(N__39151));
    InMux I__8208 (
            .O(N__39151),
            .I(N__39148));
    LocalMux I__8207 (
            .O(N__39148),
            .I(N__39145));
    Odrv12 I__8206 (
            .O(N__39145),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    InMux I__8205 (
            .O(N__39142),
            .I(N__39139));
    LocalMux I__8204 (
            .O(N__39139),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__8203 (
            .O(N__39136),
            .I(N__39133));
    LocalMux I__8202 (
            .O(N__39133),
            .I(N__39130));
    Odrv12 I__8201 (
            .O(N__39130),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__8200 (
            .O(N__39127),
            .I(N__39124));
    InMux I__8199 (
            .O(N__39124),
            .I(N__39121));
    LocalMux I__8198 (
            .O(N__39121),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__8197 (
            .O(N__39118),
            .I(N__39115));
    LocalMux I__8196 (
            .O(N__39115),
            .I(N__39112));
    Odrv12 I__8195 (
            .O(N__39112),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__8194 (
            .O(N__39109),
            .I(N__39106));
    InMux I__8193 (
            .O(N__39106),
            .I(N__39103));
    LocalMux I__8192 (
            .O(N__39103),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__8191 (
            .O(N__39100),
            .I(N__39097));
    LocalMux I__8190 (
            .O(N__39097),
            .I(N__39094));
    Odrv12 I__8189 (
            .O(N__39094),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__8188 (
            .O(N__39091),
            .I(N__39088));
    InMux I__8187 (
            .O(N__39088),
            .I(N__39085));
    LocalMux I__8186 (
            .O(N__39085),
            .I(N__39082));
    Odrv4 I__8185 (
            .O(N__39082),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    InMux I__8184 (
            .O(N__39079),
            .I(N__39076));
    LocalMux I__8183 (
            .O(N__39076),
            .I(N__39073));
    Odrv12 I__8182 (
            .O(N__39073),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__8181 (
            .O(N__39070),
            .I(N__39067));
    InMux I__8180 (
            .O(N__39067),
            .I(N__39064));
    LocalMux I__8179 (
            .O(N__39064),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__8178 (
            .O(N__39061),
            .I(N__39058));
    LocalMux I__8177 (
            .O(N__39058),
            .I(N__39055));
    Span4Mux_v I__8176 (
            .O(N__39055),
            .I(N__39052));
    Odrv4 I__8175 (
            .O(N__39052),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__8174 (
            .O(N__39049),
            .I(N__39046));
    InMux I__8173 (
            .O(N__39046),
            .I(N__39043));
    LocalMux I__8172 (
            .O(N__39043),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__8171 (
            .O(N__39040),
            .I(N__39037));
    LocalMux I__8170 (
            .O(N__39037),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__8169 (
            .O(N__39034),
            .I(N__39031));
    InMux I__8168 (
            .O(N__39031),
            .I(N__39028));
    LocalMux I__8167 (
            .O(N__39028),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__8166 (
            .O(N__39025),
            .I(N__39022));
    LocalMux I__8165 (
            .O(N__39022),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__8164 (
            .O(N__39019),
            .I(N__39016));
    InMux I__8163 (
            .O(N__39016),
            .I(N__39013));
    LocalMux I__8162 (
            .O(N__39013),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__8161 (
            .O(N__39010),
            .I(N__39007));
    LocalMux I__8160 (
            .O(N__39007),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__8159 (
            .O(N__39004),
            .I(N__39001));
    InMux I__8158 (
            .O(N__39001),
            .I(N__38998));
    LocalMux I__8157 (
            .O(N__38998),
            .I(N__38995));
    Odrv4 I__8156 (
            .O(N__38995),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__8155 (
            .O(N__38992),
            .I(N__38989));
    LocalMux I__8154 (
            .O(N__38989),
            .I(N__38986));
    Span4Mux_v I__8153 (
            .O(N__38986),
            .I(N__38983));
    Odrv4 I__8152 (
            .O(N__38983),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__8151 (
            .O(N__38980),
            .I(N__38977));
    InMux I__8150 (
            .O(N__38977),
            .I(N__38974));
    LocalMux I__8149 (
            .O(N__38974),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__8148 (
            .O(N__38971),
            .I(N__38968));
    LocalMux I__8147 (
            .O(N__38968),
            .I(N__38965));
    Span4Mux_h I__8146 (
            .O(N__38965),
            .I(N__38962));
    Odrv4 I__8145 (
            .O(N__38962),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__8144 (
            .O(N__38959),
            .I(N__38956));
    InMux I__8143 (
            .O(N__38956),
            .I(N__38953));
    LocalMux I__8142 (
            .O(N__38953),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__8141 (
            .O(N__38950),
            .I(N__38947));
    LocalMux I__8140 (
            .O(N__38947),
            .I(N__38944));
    Odrv12 I__8139 (
            .O(N__38944),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__8138 (
            .O(N__38941),
            .I(N__38938));
    InMux I__8137 (
            .O(N__38938),
            .I(N__38935));
    LocalMux I__8136 (
            .O(N__38935),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__8135 (
            .O(N__38932),
            .I(N__38929));
    LocalMux I__8134 (
            .O(N__38929),
            .I(N__38926));
    Odrv12 I__8133 (
            .O(N__38926),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__8132 (
            .O(N__38923),
            .I(N__38920));
    InMux I__8131 (
            .O(N__38920),
            .I(N__38917));
    LocalMux I__8130 (
            .O(N__38917),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    CascadeMux I__8129 (
            .O(N__38914),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_ ));
    InMux I__8128 (
            .O(N__38911),
            .I(N__38904));
    InMux I__8127 (
            .O(N__38910),
            .I(N__38904));
    InMux I__8126 (
            .O(N__38909),
            .I(N__38901));
    LocalMux I__8125 (
            .O(N__38904),
            .I(elapsed_time_ns_1_RNII6NQL1_0_1));
    LocalMux I__8124 (
            .O(N__38901),
            .I(elapsed_time_ns_1_RNII6NQL1_0_1));
    InMux I__8123 (
            .O(N__38896),
            .I(N__38892));
    InMux I__8122 (
            .O(N__38895),
            .I(N__38889));
    LocalMux I__8121 (
            .O(N__38892),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ));
    LocalMux I__8120 (
            .O(N__38889),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ));
    CascadeMux I__8119 (
            .O(N__38884),
            .I(elapsed_time_ns_1_RNII6NQL1_0_1_cascade_));
    InMux I__8118 (
            .O(N__38881),
            .I(N__38878));
    LocalMux I__8117 (
            .O(N__38878),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ));
    InMux I__8116 (
            .O(N__38875),
            .I(N__38871));
    InMux I__8115 (
            .O(N__38874),
            .I(N__38868));
    LocalMux I__8114 (
            .O(N__38871),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ));
    LocalMux I__8113 (
            .O(N__38868),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ));
    CascadeMux I__8112 (
            .O(N__38863),
            .I(elapsed_time_ns_1_RNISCJF91_0_31_cascade_));
    CascadeMux I__8111 (
            .O(N__38860),
            .I(N__38857));
    InMux I__8110 (
            .O(N__38857),
            .I(N__38852));
    CascadeMux I__8109 (
            .O(N__38856),
            .I(N__38846));
    CascadeMux I__8108 (
            .O(N__38855),
            .I(N__38840));
    LocalMux I__8107 (
            .O(N__38852),
            .I(N__38834));
    InMux I__8106 (
            .O(N__38851),
            .I(N__38829));
    InMux I__8105 (
            .O(N__38850),
            .I(N__38829));
    InMux I__8104 (
            .O(N__38849),
            .I(N__38824));
    InMux I__8103 (
            .O(N__38846),
            .I(N__38824));
    InMux I__8102 (
            .O(N__38845),
            .I(N__38819));
    InMux I__8101 (
            .O(N__38844),
            .I(N__38819));
    InMux I__8100 (
            .O(N__38843),
            .I(N__38808));
    InMux I__8099 (
            .O(N__38840),
            .I(N__38808));
    InMux I__8098 (
            .O(N__38839),
            .I(N__38808));
    InMux I__8097 (
            .O(N__38838),
            .I(N__38808));
    InMux I__8096 (
            .O(N__38837),
            .I(N__38808));
    Span4Mux_h I__8095 (
            .O(N__38834),
            .I(N__38805));
    LocalMux I__8094 (
            .O(N__38829),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__8093 (
            .O(N__38824),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__8092 (
            .O(N__38819),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    LocalMux I__8091 (
            .O(N__38808),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    Odrv4 I__8090 (
            .O(N__38805),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ));
    InMux I__8089 (
            .O(N__38794),
            .I(N__38783));
    InMux I__8088 (
            .O(N__38793),
            .I(N__38783));
    InMux I__8087 (
            .O(N__38792),
            .I(N__38783));
    CascadeMux I__8086 (
            .O(N__38791),
            .I(N__38777));
    CascadeMux I__8085 (
            .O(N__38790),
            .I(N__38773));
    LocalMux I__8084 (
            .O(N__38783),
            .I(N__38765));
    InMux I__8083 (
            .O(N__38782),
            .I(N__38760));
    InMux I__8082 (
            .O(N__38781),
            .I(N__38760));
    InMux I__8081 (
            .O(N__38780),
            .I(N__38757));
    InMux I__8080 (
            .O(N__38777),
            .I(N__38752));
    InMux I__8079 (
            .O(N__38776),
            .I(N__38752));
    InMux I__8078 (
            .O(N__38773),
            .I(N__38747));
    InMux I__8077 (
            .O(N__38772),
            .I(N__38747));
    InMux I__8076 (
            .O(N__38771),
            .I(N__38738));
    InMux I__8075 (
            .O(N__38770),
            .I(N__38738));
    InMux I__8074 (
            .O(N__38769),
            .I(N__38738));
    InMux I__8073 (
            .O(N__38768),
            .I(N__38738));
    Span4Mux_h I__8072 (
            .O(N__38765),
            .I(N__38735));
    LocalMux I__8071 (
            .O(N__38760),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__8070 (
            .O(N__38757),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__8069 (
            .O(N__38752),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__8068 (
            .O(N__38747),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    LocalMux I__8067 (
            .O(N__38738),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    Odrv4 I__8066 (
            .O(N__38735),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ));
    CascadeMux I__8065 (
            .O(N__38722),
            .I(N__38719));
    InMux I__8064 (
            .O(N__38719),
            .I(N__38716));
    LocalMux I__8063 (
            .O(N__38716),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__8062 (
            .O(N__38713),
            .I(N__38710));
    LocalMux I__8061 (
            .O(N__38710),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__8060 (
            .O(N__38707),
            .I(N__38704));
    InMux I__8059 (
            .O(N__38704),
            .I(N__38701));
    LocalMux I__8058 (
            .O(N__38701),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    InMux I__8057 (
            .O(N__38698),
            .I(N__38695));
    LocalMux I__8056 (
            .O(N__38695),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__8055 (
            .O(N__38692),
            .I(N__38689));
    LocalMux I__8054 (
            .O(N__38689),
            .I(N__38685));
    InMux I__8053 (
            .O(N__38688),
            .I(N__38680));
    Span4Mux_v I__8052 (
            .O(N__38685),
            .I(N__38677));
    InMux I__8051 (
            .O(N__38684),
            .I(N__38674));
    InMux I__8050 (
            .O(N__38683),
            .I(N__38671));
    LocalMux I__8049 (
            .O(N__38680),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ));
    Odrv4 I__8048 (
            .O(N__38677),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ));
    LocalMux I__8047 (
            .O(N__38674),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ));
    LocalMux I__8046 (
            .O(N__38671),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ));
    CascadeMux I__8045 (
            .O(N__38662),
            .I(\delay_measurement_inst.delay_tr_timer.N_386_cascade_ ));
    InMux I__8044 (
            .O(N__38659),
            .I(N__38656));
    LocalMux I__8043 (
            .O(N__38656),
            .I(N__38652));
    InMux I__8042 (
            .O(N__38655),
            .I(N__38649));
    Odrv4 I__8041 (
            .O(N__38652),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9 ));
    LocalMux I__8040 (
            .O(N__38649),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9 ));
    CascadeMux I__8039 (
            .O(N__38644),
            .I(N__38640));
    CascadeMux I__8038 (
            .O(N__38643),
            .I(N__38637));
    InMux I__8037 (
            .O(N__38640),
            .I(N__38634));
    InMux I__8036 (
            .O(N__38637),
            .I(N__38631));
    LocalMux I__8035 (
            .O(N__38634),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2 ));
    LocalMux I__8034 (
            .O(N__38631),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2 ));
    CascadeMux I__8033 (
            .O(N__38626),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2_cascade_ ));
    InMux I__8032 (
            .O(N__38623),
            .I(N__38616));
    InMux I__8031 (
            .O(N__38622),
            .I(N__38616));
    InMux I__8030 (
            .O(N__38621),
            .I(N__38613));
    LocalMux I__8029 (
            .O(N__38616),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ));
    LocalMux I__8028 (
            .O(N__38613),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ));
    InMux I__8027 (
            .O(N__38608),
            .I(N__38603));
    InMux I__8026 (
            .O(N__38607),
            .I(N__38598));
    InMux I__8025 (
            .O(N__38606),
            .I(N__38598));
    LocalMux I__8024 (
            .O(N__38603),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    LocalMux I__8023 (
            .O(N__38598),
            .I(elapsed_time_ns_1_RNIAE2591_0_2));
    InMux I__8022 (
            .O(N__38593),
            .I(N__38590));
    LocalMux I__8021 (
            .O(N__38590),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1 ));
    CascadeMux I__8020 (
            .O(N__38587),
            .I(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ));
    InMux I__8019 (
            .O(N__38584),
            .I(N__38580));
    InMux I__8018 (
            .O(N__38583),
            .I(N__38577));
    LocalMux I__8017 (
            .O(N__38580),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    LocalMux I__8016 (
            .O(N__38577),
            .I(elapsed_time_ns_1_RNI0GIF91_0_26));
    CascadeMux I__8015 (
            .O(N__38572),
            .I(N__38568));
    CascadeMux I__8014 (
            .O(N__38571),
            .I(N__38565));
    InMux I__8013 (
            .O(N__38568),
            .I(N__38561));
    InMux I__8012 (
            .O(N__38565),
            .I(N__38558));
    InMux I__8011 (
            .O(N__38564),
            .I(N__38555));
    LocalMux I__8010 (
            .O(N__38561),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    LocalMux I__8009 (
            .O(N__38558),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    LocalMux I__8008 (
            .O(N__38555),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10));
    InMux I__8007 (
            .O(N__38548),
            .I(N__38542));
    InMux I__8006 (
            .O(N__38547),
            .I(N__38539));
    InMux I__8005 (
            .O(N__38546),
            .I(N__38536));
    InMux I__8004 (
            .O(N__38545),
            .I(N__38533));
    LocalMux I__8003 (
            .O(N__38542),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    LocalMux I__8002 (
            .O(N__38539),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    LocalMux I__8001 (
            .O(N__38536),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    LocalMux I__8000 (
            .O(N__38533),
            .I(elapsed_time_ns_1_RNIQ8HF91_0_11));
    InMux I__7999 (
            .O(N__38524),
            .I(N__38518));
    InMux I__7998 (
            .O(N__38523),
            .I(N__38515));
    InMux I__7997 (
            .O(N__38522),
            .I(N__38512));
    InMux I__7996 (
            .O(N__38521),
            .I(N__38509));
    LocalMux I__7995 (
            .O(N__38518),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__7994 (
            .O(N__38515),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__7993 (
            .O(N__38512),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    LocalMux I__7992 (
            .O(N__38509),
            .I(elapsed_time_ns_1_RNIR9HF91_0_12));
    CascadeMux I__7991 (
            .O(N__38500),
            .I(N__38496));
    InMux I__7990 (
            .O(N__38499),
            .I(N__38491));
    InMux I__7989 (
            .O(N__38496),
            .I(N__38488));
    InMux I__7988 (
            .O(N__38495),
            .I(N__38485));
    InMux I__7987 (
            .O(N__38494),
            .I(N__38482));
    LocalMux I__7986 (
            .O(N__38491),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    LocalMux I__7985 (
            .O(N__38488),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    LocalMux I__7984 (
            .O(N__38485),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    LocalMux I__7983 (
            .O(N__38482),
            .I(elapsed_time_ns_1_RNISAHF91_0_13));
    InMux I__7982 (
            .O(N__38473),
            .I(N__38462));
    InMux I__7981 (
            .O(N__38472),
            .I(N__38462));
    InMux I__7980 (
            .O(N__38471),
            .I(N__38459));
    InMux I__7979 (
            .O(N__38470),
            .I(N__38456));
    InMux I__7978 (
            .O(N__38469),
            .I(N__38453));
    InMux I__7977 (
            .O(N__38468),
            .I(N__38448));
    InMux I__7976 (
            .O(N__38467),
            .I(N__38448));
    LocalMux I__7975 (
            .O(N__38462),
            .I(N__38445));
    LocalMux I__7974 (
            .O(N__38459),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__7973 (
            .O(N__38456),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__7972 (
            .O(N__38453),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    LocalMux I__7971 (
            .O(N__38448),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    Odrv4 I__7970 (
            .O(N__38445),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15));
    CascadeMux I__7969 (
            .O(N__38434),
            .I(elapsed_time_ns_1_RNIUCHF91_0_15_cascade_));
    CascadeMux I__7968 (
            .O(N__38431),
            .I(N__38423));
    CascadeMux I__7967 (
            .O(N__38430),
            .I(N__38420));
    InMux I__7966 (
            .O(N__38429),
            .I(N__38411));
    InMux I__7965 (
            .O(N__38428),
            .I(N__38400));
    InMux I__7964 (
            .O(N__38427),
            .I(N__38400));
    InMux I__7963 (
            .O(N__38426),
            .I(N__38400));
    InMux I__7962 (
            .O(N__38423),
            .I(N__38400));
    InMux I__7961 (
            .O(N__38420),
            .I(N__38400));
    InMux I__7960 (
            .O(N__38419),
            .I(N__38387));
    InMux I__7959 (
            .O(N__38418),
            .I(N__38387));
    InMux I__7958 (
            .O(N__38417),
            .I(N__38387));
    InMux I__7957 (
            .O(N__38416),
            .I(N__38387));
    InMux I__7956 (
            .O(N__38415),
            .I(N__38387));
    InMux I__7955 (
            .O(N__38414),
            .I(N__38387));
    LocalMux I__7954 (
            .O(N__38411),
            .I(\phase_controller_inst1.stoper_tr.N_244 ));
    LocalMux I__7953 (
            .O(N__38400),
            .I(\phase_controller_inst1.stoper_tr.N_244 ));
    LocalMux I__7952 (
            .O(N__38387),
            .I(\phase_controller_inst1.stoper_tr.N_244 ));
    InMux I__7951 (
            .O(N__38380),
            .I(N__38377));
    LocalMux I__7950 (
            .O(N__38377),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ));
    InMux I__7949 (
            .O(N__38374),
            .I(N__38371));
    LocalMux I__7948 (
            .O(N__38371),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25));
    CascadeMux I__7947 (
            .O(N__38368),
            .I(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_));
    InMux I__7946 (
            .O(N__38365),
            .I(N__38359));
    InMux I__7945 (
            .O(N__38364),
            .I(N__38359));
    LocalMux I__7944 (
            .O(N__38359),
            .I(elapsed_time_ns_1_RNI2IIF91_0_28));
    CascadeMux I__7943 (
            .O(N__38356),
            .I(N__38353));
    InMux I__7942 (
            .O(N__38353),
            .I(N__38347));
    InMux I__7941 (
            .O(N__38352),
            .I(N__38347));
    LocalMux I__7940 (
            .O(N__38347),
            .I(elapsed_time_ns_1_RNI1HIF91_0_27));
    InMux I__7939 (
            .O(N__38344),
            .I(N__38341));
    LocalMux I__7938 (
            .O(N__38341),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15 ));
    CascadeMux I__7937 (
            .O(N__38338),
            .I(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_ ));
    CascadeMux I__7936 (
            .O(N__38335),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ));
    InMux I__7935 (
            .O(N__38332),
            .I(N__38326));
    InMux I__7934 (
            .O(N__38331),
            .I(N__38326));
    LocalMux I__7933 (
            .O(N__38326),
            .I(elapsed_time_ns_1_RNISBIF91_0_22));
    CascadeMux I__7932 (
            .O(N__38323),
            .I(N__38319));
    InMux I__7931 (
            .O(N__38322),
            .I(N__38316));
    InMux I__7930 (
            .O(N__38319),
            .I(N__38313));
    LocalMux I__7929 (
            .O(N__38316),
            .I(N__38309));
    LocalMux I__7928 (
            .O(N__38313),
            .I(N__38306));
    InMux I__7927 (
            .O(N__38312),
            .I(N__38303));
    Odrv4 I__7926 (
            .O(N__38309),
            .I(elapsed_time_ns_1_RNIOJKEE1_0_7));
    Odrv4 I__7925 (
            .O(N__38306),
            .I(elapsed_time_ns_1_RNIOJKEE1_0_7));
    LocalMux I__7924 (
            .O(N__38303),
            .I(elapsed_time_ns_1_RNIOJKEE1_0_7));
    CascadeMux I__7923 (
            .O(N__38296),
            .I(N__38291));
    InMux I__7922 (
            .O(N__38295),
            .I(N__38288));
    InMux I__7921 (
            .O(N__38294),
            .I(N__38285));
    InMux I__7920 (
            .O(N__38291),
            .I(N__38282));
    LocalMux I__7919 (
            .O(N__38288),
            .I(N__38279));
    LocalMux I__7918 (
            .O(N__38285),
            .I(N__38274));
    LocalMux I__7917 (
            .O(N__38282),
            .I(N__38274));
    Span4Mux_h I__7916 (
            .O(N__38279),
            .I(N__38271));
    Span12Mux_h I__7915 (
            .O(N__38274),
            .I(N__38266));
    Sp12to4 I__7914 (
            .O(N__38271),
            .I(N__38266));
    Span12Mux_v I__7913 (
            .O(N__38266),
            .I(N__38263));
    Odrv12 I__7912 (
            .O(N__38263),
            .I(il_max_comp1_D2));
    InMux I__7911 (
            .O(N__38260),
            .I(N__38247));
    InMux I__7910 (
            .O(N__38259),
            .I(N__38247));
    InMux I__7909 (
            .O(N__38258),
            .I(N__38247));
    InMux I__7908 (
            .O(N__38257),
            .I(N__38243));
    InMux I__7907 (
            .O(N__38256),
            .I(N__38240));
    InMux I__7906 (
            .O(N__38255),
            .I(N__38237));
    InMux I__7905 (
            .O(N__38254),
            .I(N__38234));
    LocalMux I__7904 (
            .O(N__38247),
            .I(N__38231));
    InMux I__7903 (
            .O(N__38246),
            .I(N__38228));
    LocalMux I__7902 (
            .O(N__38243),
            .I(state_3));
    LocalMux I__7901 (
            .O(N__38240),
            .I(state_3));
    LocalMux I__7900 (
            .O(N__38237),
            .I(state_3));
    LocalMux I__7899 (
            .O(N__38234),
            .I(state_3));
    Odrv4 I__7898 (
            .O(N__38231),
            .I(state_3));
    LocalMux I__7897 (
            .O(N__38228),
            .I(state_3));
    IoInMux I__7896 (
            .O(N__38215),
            .I(N__38212));
    LocalMux I__7895 (
            .O(N__38212),
            .I(N__38209));
    IoSpan4Mux I__7894 (
            .O(N__38209),
            .I(N__38206));
    Span4Mux_s3_v I__7893 (
            .O(N__38206),
            .I(N__38203));
    Span4Mux_v I__7892 (
            .O(N__38203),
            .I(N__38199));
    InMux I__7891 (
            .O(N__38202),
            .I(N__38196));
    Odrv4 I__7890 (
            .O(N__38199),
            .I(T01_c));
    LocalMux I__7889 (
            .O(N__38196),
            .I(T01_c));
    InMux I__7888 (
            .O(N__38191),
            .I(N__38188));
    LocalMux I__7887 (
            .O(N__38188),
            .I(N__38185));
    Span4Mux_h I__7886 (
            .O(N__38185),
            .I(N__38182));
    Odrv4 I__7885 (
            .O(N__38182),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    CascadeMux I__7884 (
            .O(N__38179),
            .I(N__38175));
    CascadeMux I__7883 (
            .O(N__38178),
            .I(N__38171));
    InMux I__7882 (
            .O(N__38175),
            .I(N__38168));
    CascadeMux I__7881 (
            .O(N__38174),
            .I(N__38165));
    InMux I__7880 (
            .O(N__38171),
            .I(N__38162));
    LocalMux I__7879 (
            .O(N__38168),
            .I(N__38159));
    InMux I__7878 (
            .O(N__38165),
            .I(N__38156));
    LocalMux I__7877 (
            .O(N__38162),
            .I(N__38151));
    Span4Mux_v I__7876 (
            .O(N__38159),
            .I(N__38146));
    LocalMux I__7875 (
            .O(N__38156),
            .I(N__38146));
    InMux I__7874 (
            .O(N__38155),
            .I(N__38141));
    InMux I__7873 (
            .O(N__38154),
            .I(N__38141));
    Span4Mux_h I__7872 (
            .O(N__38151),
            .I(N__38138));
    Span4Mux_h I__7871 (
            .O(N__38146),
            .I(N__38133));
    LocalMux I__7870 (
            .O(N__38141),
            .I(N__38133));
    Span4Mux_h I__7869 (
            .O(N__38138),
            .I(N__38130));
    Span4Mux_h I__7868 (
            .O(N__38133),
            .I(N__38127));
    Odrv4 I__7867 (
            .O(N__38130),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__7866 (
            .O(N__38127),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__7865 (
            .O(N__38122),
            .I(N__38119));
    LocalMux I__7864 (
            .O(N__38119),
            .I(N__38116));
    Span4Mux_h I__7863 (
            .O(N__38116),
            .I(N__38113));
    Odrv4 I__7862 (
            .O(N__38113),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    CascadeMux I__7861 (
            .O(N__38110),
            .I(N__38107));
    InMux I__7860 (
            .O(N__38107),
            .I(N__38104));
    LocalMux I__7859 (
            .O(N__38104),
            .I(N__38100));
    InMux I__7858 (
            .O(N__38103),
            .I(N__38097));
    Span4Mux_h I__7857 (
            .O(N__38100),
            .I(N__38090));
    LocalMux I__7856 (
            .O(N__38097),
            .I(N__38090));
    InMux I__7855 (
            .O(N__38096),
            .I(N__38087));
    InMux I__7854 (
            .O(N__38095),
            .I(N__38083));
    Span4Mux_v I__7853 (
            .O(N__38090),
            .I(N__38080));
    LocalMux I__7852 (
            .O(N__38087),
            .I(N__38077));
    InMux I__7851 (
            .O(N__38086),
            .I(N__38074));
    LocalMux I__7850 (
            .O(N__38083),
            .I(N__38069));
    Sp12to4 I__7849 (
            .O(N__38080),
            .I(N__38069));
    Span4Mux_h I__7848 (
            .O(N__38077),
            .I(N__38064));
    LocalMux I__7847 (
            .O(N__38074),
            .I(N__38064));
    Odrv12 I__7846 (
            .O(N__38069),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__7845 (
            .O(N__38064),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__7844 (
            .O(N__38059),
            .I(N__38054));
    InMux I__7843 (
            .O(N__38058),
            .I(N__38051));
    InMux I__7842 (
            .O(N__38057),
            .I(N__38048));
    LocalMux I__7841 (
            .O(N__38054),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    LocalMux I__7840 (
            .O(N__38051),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    LocalMux I__7839 (
            .O(N__38048),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ));
    CascadeMux I__7838 (
            .O(N__38041),
            .I(N__38038));
    InMux I__7837 (
            .O(N__38038),
            .I(N__38032));
    InMux I__7836 (
            .O(N__38037),
            .I(N__38029));
    InMux I__7835 (
            .O(N__38036),
            .I(N__38026));
    InMux I__7834 (
            .O(N__38035),
            .I(N__38023));
    LocalMux I__7833 (
            .O(N__38032),
            .I(N__38020));
    LocalMux I__7832 (
            .O(N__38029),
            .I(N__38017));
    LocalMux I__7831 (
            .O(N__38026),
            .I(N__38014));
    LocalMux I__7830 (
            .O(N__38023),
            .I(N__38011));
    Span4Mux_v I__7829 (
            .O(N__38020),
            .I(N__38008));
    Span4Mux_v I__7828 (
            .O(N__38017),
            .I(N__38005));
    Span4Mux_h I__7827 (
            .O(N__38014),
            .I(N__38001));
    Span4Mux_v I__7826 (
            .O(N__38011),
            .I(N__37994));
    Span4Mux_h I__7825 (
            .O(N__38008),
            .I(N__37994));
    Span4Mux_h I__7824 (
            .O(N__38005),
            .I(N__37994));
    InMux I__7823 (
            .O(N__38004),
            .I(N__37991));
    Odrv4 I__7822 (
            .O(N__38001),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv4 I__7821 (
            .O(N__37994),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__7820 (
            .O(N__37991),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    CascadeMux I__7819 (
            .O(N__37984),
            .I(N__37980));
    InMux I__7818 (
            .O(N__37983),
            .I(N__37966));
    InMux I__7817 (
            .O(N__37980),
            .I(N__37963));
    InMux I__7816 (
            .O(N__37979),
            .I(N__37954));
    InMux I__7815 (
            .O(N__37978),
            .I(N__37954));
    InMux I__7814 (
            .O(N__37977),
            .I(N__37954));
    InMux I__7813 (
            .O(N__37976),
            .I(N__37954));
    CascadeMux I__7812 (
            .O(N__37975),
            .I(N__37951));
    InMux I__7811 (
            .O(N__37974),
            .I(N__37919));
    InMux I__7810 (
            .O(N__37973),
            .I(N__37919));
    InMux I__7809 (
            .O(N__37972),
            .I(N__37919));
    InMux I__7808 (
            .O(N__37971),
            .I(N__37919));
    InMux I__7807 (
            .O(N__37970),
            .I(N__37919));
    InMux I__7806 (
            .O(N__37969),
            .I(N__37919));
    LocalMux I__7805 (
            .O(N__37966),
            .I(N__37916));
    LocalMux I__7804 (
            .O(N__37963),
            .I(N__37911));
    LocalMux I__7803 (
            .O(N__37954),
            .I(N__37911));
    InMux I__7802 (
            .O(N__37951),
            .I(N__37900));
    InMux I__7801 (
            .O(N__37950),
            .I(N__37900));
    InMux I__7800 (
            .O(N__37949),
            .I(N__37900));
    InMux I__7799 (
            .O(N__37948),
            .I(N__37900));
    InMux I__7798 (
            .O(N__37947),
            .I(N__37900));
    InMux I__7797 (
            .O(N__37946),
            .I(N__37897));
    CascadeMux I__7796 (
            .O(N__37945),
            .I(N__37894));
    CascadeMux I__7795 (
            .O(N__37944),
            .I(N__37889));
    CascadeMux I__7794 (
            .O(N__37943),
            .I(N__37885));
    CascadeMux I__7793 (
            .O(N__37942),
            .I(N__37879));
    CascadeMux I__7792 (
            .O(N__37941),
            .I(N__37874));
    CascadeMux I__7791 (
            .O(N__37940),
            .I(N__37868));
    InMux I__7790 (
            .O(N__37939),
            .I(N__37860));
    InMux I__7789 (
            .O(N__37938),
            .I(N__37860));
    InMux I__7788 (
            .O(N__37937),
            .I(N__37860));
    InMux I__7787 (
            .O(N__37936),
            .I(N__37851));
    InMux I__7786 (
            .O(N__37935),
            .I(N__37851));
    InMux I__7785 (
            .O(N__37934),
            .I(N__37851));
    InMux I__7784 (
            .O(N__37933),
            .I(N__37851));
    InMux I__7783 (
            .O(N__37932),
            .I(N__37848));
    LocalMux I__7782 (
            .O(N__37919),
            .I(N__37839));
    Span4Mux_v I__7781 (
            .O(N__37916),
            .I(N__37839));
    Span4Mux_v I__7780 (
            .O(N__37911),
            .I(N__37839));
    LocalMux I__7779 (
            .O(N__37900),
            .I(N__37839));
    LocalMux I__7778 (
            .O(N__37897),
            .I(N__37834));
    InMux I__7777 (
            .O(N__37894),
            .I(N__37828));
    InMux I__7776 (
            .O(N__37893),
            .I(N__37828));
    InMux I__7775 (
            .O(N__37892),
            .I(N__37817));
    InMux I__7774 (
            .O(N__37889),
            .I(N__37817));
    InMux I__7773 (
            .O(N__37888),
            .I(N__37817));
    InMux I__7772 (
            .O(N__37885),
            .I(N__37817));
    InMux I__7771 (
            .O(N__37884),
            .I(N__37817));
    InMux I__7770 (
            .O(N__37883),
            .I(N__37806));
    InMux I__7769 (
            .O(N__37882),
            .I(N__37806));
    InMux I__7768 (
            .O(N__37879),
            .I(N__37806));
    InMux I__7767 (
            .O(N__37878),
            .I(N__37806));
    InMux I__7766 (
            .O(N__37877),
            .I(N__37806));
    InMux I__7765 (
            .O(N__37874),
            .I(N__37793));
    InMux I__7764 (
            .O(N__37873),
            .I(N__37793));
    InMux I__7763 (
            .O(N__37872),
            .I(N__37793));
    InMux I__7762 (
            .O(N__37871),
            .I(N__37793));
    InMux I__7761 (
            .O(N__37868),
            .I(N__37793));
    InMux I__7760 (
            .O(N__37867),
            .I(N__37793));
    LocalMux I__7759 (
            .O(N__37860),
            .I(N__37786));
    LocalMux I__7758 (
            .O(N__37851),
            .I(N__37786));
    LocalMux I__7757 (
            .O(N__37848),
            .I(N__37781));
    Span4Mux_h I__7756 (
            .O(N__37839),
            .I(N__37781));
    InMux I__7755 (
            .O(N__37838),
            .I(N__37776));
    InMux I__7754 (
            .O(N__37837),
            .I(N__37776));
    Span4Mux_h I__7753 (
            .O(N__37834),
            .I(N__37773));
    InMux I__7752 (
            .O(N__37833),
            .I(N__37770));
    LocalMux I__7751 (
            .O(N__37828),
            .I(N__37761));
    LocalMux I__7750 (
            .O(N__37817),
            .I(N__37761));
    LocalMux I__7749 (
            .O(N__37806),
            .I(N__37761));
    LocalMux I__7748 (
            .O(N__37793),
            .I(N__37761));
    InMux I__7747 (
            .O(N__37792),
            .I(N__37756));
    InMux I__7746 (
            .O(N__37791),
            .I(N__37756));
    Span4Mux_v I__7745 (
            .O(N__37786),
            .I(N__37751));
    Span4Mux_v I__7744 (
            .O(N__37781),
            .I(N__37751));
    LocalMux I__7743 (
            .O(N__37776),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__7742 (
            .O(N__37773),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    LocalMux I__7741 (
            .O(N__37770),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv12 I__7740 (
            .O(N__37761),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    LocalMux I__7739 (
            .O(N__37756),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv4 I__7738 (
            .O(N__37751),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__7737 (
            .O(N__37738),
            .I(N__37735));
    LocalMux I__7736 (
            .O(N__37735),
            .I(N__37732));
    Odrv4 I__7735 (
            .O(N__37732),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ));
    CascadeMux I__7734 (
            .O(N__37729),
            .I(N__37726));
    InMux I__7733 (
            .O(N__37726),
            .I(N__37723));
    LocalMux I__7732 (
            .O(N__37723),
            .I(N__37720));
    Span4Mux_h I__7731 (
            .O(N__37720),
            .I(N__37717));
    Odrv4 I__7730 (
            .O(N__37717),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0 ));
    CascadeMux I__7729 (
            .O(N__37714),
            .I(N__37710));
    InMux I__7728 (
            .O(N__37713),
            .I(N__37703));
    InMux I__7727 (
            .O(N__37710),
            .I(N__37700));
    InMux I__7726 (
            .O(N__37709),
            .I(N__37697));
    CascadeMux I__7725 (
            .O(N__37708),
            .I(N__37694));
    InMux I__7724 (
            .O(N__37707),
            .I(N__37689));
    CascadeMux I__7723 (
            .O(N__37706),
            .I(N__37683));
    LocalMux I__7722 (
            .O(N__37703),
            .I(N__37674));
    LocalMux I__7721 (
            .O(N__37700),
            .I(N__37674));
    LocalMux I__7720 (
            .O(N__37697),
            .I(N__37674));
    InMux I__7719 (
            .O(N__37694),
            .I(N__37660));
    InMux I__7718 (
            .O(N__37693),
            .I(N__37655));
    InMux I__7717 (
            .O(N__37692),
            .I(N__37655));
    LocalMux I__7716 (
            .O(N__37689),
            .I(N__37652));
    InMux I__7715 (
            .O(N__37688),
            .I(N__37643));
    InMux I__7714 (
            .O(N__37687),
            .I(N__37643));
    InMux I__7713 (
            .O(N__37686),
            .I(N__37643));
    InMux I__7712 (
            .O(N__37683),
            .I(N__37643));
    InMux I__7711 (
            .O(N__37682),
            .I(N__37640));
    InMux I__7710 (
            .O(N__37681),
            .I(N__37637));
    Span4Mux_v I__7709 (
            .O(N__37674),
            .I(N__37634));
    InMux I__7708 (
            .O(N__37673),
            .I(N__37631));
    CascadeMux I__7707 (
            .O(N__37672),
            .I(N__37624));
    CascadeMux I__7706 (
            .O(N__37671),
            .I(N__37621));
    CascadeMux I__7705 (
            .O(N__37670),
            .I(N__37618));
    CascadeMux I__7704 (
            .O(N__37669),
            .I(N__37615));
    CascadeMux I__7703 (
            .O(N__37668),
            .I(N__37609));
    CascadeMux I__7702 (
            .O(N__37667),
            .I(N__37606));
    InMux I__7701 (
            .O(N__37666),
            .I(N__37603));
    CascadeMux I__7700 (
            .O(N__37665),
            .I(N__37599));
    InMux I__7699 (
            .O(N__37664),
            .I(N__37596));
    InMux I__7698 (
            .O(N__37663),
            .I(N__37593));
    LocalMux I__7697 (
            .O(N__37660),
            .I(N__37588));
    LocalMux I__7696 (
            .O(N__37655),
            .I(N__37588));
    Span4Mux_v I__7695 (
            .O(N__37652),
            .I(N__37583));
    LocalMux I__7694 (
            .O(N__37643),
            .I(N__37583));
    LocalMux I__7693 (
            .O(N__37640),
            .I(N__37578));
    LocalMux I__7692 (
            .O(N__37637),
            .I(N__37578));
    Span4Mux_h I__7691 (
            .O(N__37634),
            .I(N__37573));
    LocalMux I__7690 (
            .O(N__37631),
            .I(N__37573));
    InMux I__7689 (
            .O(N__37630),
            .I(N__37556));
    InMux I__7688 (
            .O(N__37629),
            .I(N__37556));
    InMux I__7687 (
            .O(N__37628),
            .I(N__37556));
    InMux I__7686 (
            .O(N__37627),
            .I(N__37556));
    InMux I__7685 (
            .O(N__37624),
            .I(N__37556));
    InMux I__7684 (
            .O(N__37621),
            .I(N__37556));
    InMux I__7683 (
            .O(N__37618),
            .I(N__37556));
    InMux I__7682 (
            .O(N__37615),
            .I(N__37556));
    InMux I__7681 (
            .O(N__37614),
            .I(N__37545));
    InMux I__7680 (
            .O(N__37613),
            .I(N__37545));
    InMux I__7679 (
            .O(N__37612),
            .I(N__37545));
    InMux I__7678 (
            .O(N__37609),
            .I(N__37545));
    InMux I__7677 (
            .O(N__37606),
            .I(N__37545));
    LocalMux I__7676 (
            .O(N__37603),
            .I(N__37542));
    InMux I__7675 (
            .O(N__37602),
            .I(N__37537));
    InMux I__7674 (
            .O(N__37599),
            .I(N__37537));
    LocalMux I__7673 (
            .O(N__37596),
            .I(N__37530));
    LocalMux I__7672 (
            .O(N__37593),
            .I(N__37530));
    Span4Mux_h I__7671 (
            .O(N__37588),
            .I(N__37530));
    Span4Mux_h I__7670 (
            .O(N__37583),
            .I(N__37527));
    Span12Mux_h I__7669 (
            .O(N__37578),
            .I(N__37524));
    Span4Mux_h I__7668 (
            .O(N__37573),
            .I(N__37521));
    LocalMux I__7667 (
            .O(N__37556),
            .I(N__37514));
    LocalMux I__7666 (
            .O(N__37545),
            .I(N__37514));
    Span12Mux_s7_v I__7665 (
            .O(N__37542),
            .I(N__37514));
    LocalMux I__7664 (
            .O(N__37537),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__7663 (
            .O(N__37530),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__7662 (
            .O(N__37527),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv12 I__7661 (
            .O(N__37524),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv4 I__7660 (
            .O(N__37521),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    Odrv12 I__7659 (
            .O(N__37514),
            .I(\current_shift_inst.PI_CTRL.N_74 ));
    InMux I__7658 (
            .O(N__37501),
            .I(N__37489));
    InMux I__7657 (
            .O(N__37500),
            .I(N__37485));
    InMux I__7656 (
            .O(N__37499),
            .I(N__37482));
    InMux I__7655 (
            .O(N__37498),
            .I(N__37479));
    InMux I__7654 (
            .O(N__37497),
            .I(N__37476));
    InMux I__7653 (
            .O(N__37496),
            .I(N__37464));
    InMux I__7652 (
            .O(N__37495),
            .I(N__37464));
    InMux I__7651 (
            .O(N__37494),
            .I(N__37464));
    InMux I__7650 (
            .O(N__37493),
            .I(N__37464));
    InMux I__7649 (
            .O(N__37492),
            .I(N__37464));
    LocalMux I__7648 (
            .O(N__37489),
            .I(N__37461));
    InMux I__7647 (
            .O(N__37488),
            .I(N__37457));
    LocalMux I__7646 (
            .O(N__37485),
            .I(N__37435));
    LocalMux I__7645 (
            .O(N__37482),
            .I(N__37432));
    LocalMux I__7644 (
            .O(N__37479),
            .I(N__37427));
    LocalMux I__7643 (
            .O(N__37476),
            .I(N__37427));
    InMux I__7642 (
            .O(N__37475),
            .I(N__37424));
    LocalMux I__7641 (
            .O(N__37464),
            .I(N__37419));
    Span4Mux_h I__7640 (
            .O(N__37461),
            .I(N__37419));
    InMux I__7639 (
            .O(N__37460),
            .I(N__37416));
    LocalMux I__7638 (
            .O(N__37457),
            .I(N__37413));
    InMux I__7637 (
            .O(N__37456),
            .I(N__37404));
    InMux I__7636 (
            .O(N__37455),
            .I(N__37404));
    InMux I__7635 (
            .O(N__37454),
            .I(N__37404));
    InMux I__7634 (
            .O(N__37453),
            .I(N__37404));
    InMux I__7633 (
            .O(N__37452),
            .I(N__37387));
    InMux I__7632 (
            .O(N__37451),
            .I(N__37387));
    InMux I__7631 (
            .O(N__37450),
            .I(N__37387));
    InMux I__7630 (
            .O(N__37449),
            .I(N__37387));
    InMux I__7629 (
            .O(N__37448),
            .I(N__37387));
    InMux I__7628 (
            .O(N__37447),
            .I(N__37387));
    InMux I__7627 (
            .O(N__37446),
            .I(N__37387));
    InMux I__7626 (
            .O(N__37445),
            .I(N__37387));
    InMux I__7625 (
            .O(N__37444),
            .I(N__37384));
    InMux I__7624 (
            .O(N__37443),
            .I(N__37377));
    InMux I__7623 (
            .O(N__37442),
            .I(N__37377));
    InMux I__7622 (
            .O(N__37441),
            .I(N__37377));
    InMux I__7621 (
            .O(N__37440),
            .I(N__37372));
    InMux I__7620 (
            .O(N__37439),
            .I(N__37372));
    InMux I__7619 (
            .O(N__37438),
            .I(N__37369));
    Span4Mux_v I__7618 (
            .O(N__37435),
            .I(N__37366));
    Span4Mux_v I__7617 (
            .O(N__37432),
            .I(N__37363));
    Span12Mux_s9_v I__7616 (
            .O(N__37427),
            .I(N__37360));
    LocalMux I__7615 (
            .O(N__37424),
            .I(N__37351));
    Span4Mux_v I__7614 (
            .O(N__37419),
            .I(N__37351));
    LocalMux I__7613 (
            .O(N__37416),
            .I(N__37351));
    Span4Mux_v I__7612 (
            .O(N__37413),
            .I(N__37351));
    LocalMux I__7611 (
            .O(N__37404),
            .I(N__37344));
    LocalMux I__7610 (
            .O(N__37387),
            .I(N__37344));
    LocalMux I__7609 (
            .O(N__37384),
            .I(N__37344));
    LocalMux I__7608 (
            .O(N__37377),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__7607 (
            .O(N__37372),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__7606 (
            .O(N__37369),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__7605 (
            .O(N__37366),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__7604 (
            .O(N__37363),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__7603 (
            .O(N__37360),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__7602 (
            .O(N__37351),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__7601 (
            .O(N__37344),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    CascadeMux I__7600 (
            .O(N__37327),
            .I(N__37320));
    CascadeMux I__7599 (
            .O(N__37326),
            .I(N__37317));
    CascadeMux I__7598 (
            .O(N__37325),
            .I(N__37312));
    CascadeMux I__7597 (
            .O(N__37324),
            .I(N__37309));
    InMux I__7596 (
            .O(N__37323),
            .I(N__37304));
    InMux I__7595 (
            .O(N__37320),
            .I(N__37300));
    InMux I__7594 (
            .O(N__37317),
            .I(N__37297));
    InMux I__7593 (
            .O(N__37316),
            .I(N__37294));
    InMux I__7592 (
            .O(N__37315),
            .I(N__37291));
    InMux I__7591 (
            .O(N__37312),
            .I(N__37277));
    InMux I__7590 (
            .O(N__37309),
            .I(N__37277));
    InMux I__7589 (
            .O(N__37308),
            .I(N__37274));
    InMux I__7588 (
            .O(N__37307),
            .I(N__37263));
    LocalMux I__7587 (
            .O(N__37304),
            .I(N__37260));
    InMux I__7586 (
            .O(N__37303),
            .I(N__37257));
    LocalMux I__7585 (
            .O(N__37300),
            .I(N__37254));
    LocalMux I__7584 (
            .O(N__37297),
            .I(N__37251));
    LocalMux I__7583 (
            .O(N__37294),
            .I(N__37246));
    LocalMux I__7582 (
            .O(N__37291),
            .I(N__37246));
    InMux I__7581 (
            .O(N__37290),
            .I(N__37235));
    InMux I__7580 (
            .O(N__37289),
            .I(N__37235));
    InMux I__7579 (
            .O(N__37288),
            .I(N__37235));
    InMux I__7578 (
            .O(N__37287),
            .I(N__37235));
    InMux I__7577 (
            .O(N__37286),
            .I(N__37235));
    InMux I__7576 (
            .O(N__37285),
            .I(N__37227));
    InMux I__7575 (
            .O(N__37284),
            .I(N__37224));
    InMux I__7574 (
            .O(N__37283),
            .I(N__37219));
    InMux I__7573 (
            .O(N__37282),
            .I(N__37219));
    LocalMux I__7572 (
            .O(N__37277),
            .I(N__37216));
    LocalMux I__7571 (
            .O(N__37274),
            .I(N__37213));
    InMux I__7570 (
            .O(N__37273),
            .I(N__37196));
    InMux I__7569 (
            .O(N__37272),
            .I(N__37196));
    InMux I__7568 (
            .O(N__37271),
            .I(N__37196));
    InMux I__7567 (
            .O(N__37270),
            .I(N__37196));
    InMux I__7566 (
            .O(N__37269),
            .I(N__37196));
    InMux I__7565 (
            .O(N__37268),
            .I(N__37196));
    InMux I__7564 (
            .O(N__37267),
            .I(N__37196));
    InMux I__7563 (
            .O(N__37266),
            .I(N__37196));
    LocalMux I__7562 (
            .O(N__37263),
            .I(N__37191));
    Span4Mux_h I__7561 (
            .O(N__37260),
            .I(N__37191));
    LocalMux I__7560 (
            .O(N__37257),
            .I(N__37188));
    Span4Mux_v I__7559 (
            .O(N__37254),
            .I(N__37183));
    Span4Mux_v I__7558 (
            .O(N__37251),
            .I(N__37183));
    Span4Mux_h I__7557 (
            .O(N__37246),
            .I(N__37178));
    LocalMux I__7556 (
            .O(N__37235),
            .I(N__37178));
    InMux I__7555 (
            .O(N__37234),
            .I(N__37175));
    InMux I__7554 (
            .O(N__37233),
            .I(N__37166));
    InMux I__7553 (
            .O(N__37232),
            .I(N__37166));
    InMux I__7552 (
            .O(N__37231),
            .I(N__37166));
    InMux I__7551 (
            .O(N__37230),
            .I(N__37166));
    LocalMux I__7550 (
            .O(N__37227),
            .I(N__37161));
    LocalMux I__7549 (
            .O(N__37224),
            .I(N__37161));
    LocalMux I__7548 (
            .O(N__37219),
            .I(N__37158));
    Span4Mux_v I__7547 (
            .O(N__37216),
            .I(N__37151));
    Span4Mux_v I__7546 (
            .O(N__37213),
            .I(N__37151));
    LocalMux I__7545 (
            .O(N__37196),
            .I(N__37151));
    Span4Mux_h I__7544 (
            .O(N__37191),
            .I(N__37148));
    Span4Mux_v I__7543 (
            .O(N__37188),
            .I(N__37143));
    Span4Mux_h I__7542 (
            .O(N__37183),
            .I(N__37143));
    Span4Mux_v I__7541 (
            .O(N__37178),
            .I(N__37140));
    LocalMux I__7540 (
            .O(N__37175),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    LocalMux I__7539 (
            .O(N__37166),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv12 I__7538 (
            .O(N__37161),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv12 I__7537 (
            .O(N__37158),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__7536 (
            .O(N__37151),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__7535 (
            .O(N__37148),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__7534 (
            .O(N__37143),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    Odrv4 I__7533 (
            .O(N__37140),
            .I(\current_shift_inst.PI_CTRL.N_75 ));
    InMux I__7532 (
            .O(N__37123),
            .I(N__37120));
    LocalMux I__7531 (
            .O(N__37120),
            .I(N__37117));
    Odrv12 I__7530 (
            .O(N__37117),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    CascadeMux I__7529 (
            .O(N__37114),
            .I(N__37111));
    InMux I__7528 (
            .O(N__37111),
            .I(N__37108));
    LocalMux I__7527 (
            .O(N__37108),
            .I(N__37104));
    InMux I__7526 (
            .O(N__37107),
            .I(N__37101));
    Span4Mux_h I__7525 (
            .O(N__37104),
            .I(N__37095));
    LocalMux I__7524 (
            .O(N__37101),
            .I(N__37095));
    InMux I__7523 (
            .O(N__37100),
            .I(N__37092));
    Span4Mux_v I__7522 (
            .O(N__37095),
            .I(N__37086));
    LocalMux I__7521 (
            .O(N__37092),
            .I(N__37086));
    InMux I__7520 (
            .O(N__37091),
            .I(N__37083));
    Span4Mux_h I__7519 (
            .O(N__37086),
            .I(N__37079));
    LocalMux I__7518 (
            .O(N__37083),
            .I(N__37076));
    InMux I__7517 (
            .O(N__37082),
            .I(N__37073));
    Span4Mux_h I__7516 (
            .O(N__37079),
            .I(N__37070));
    Span4Mux_h I__7515 (
            .O(N__37076),
            .I(N__37067));
    LocalMux I__7514 (
            .O(N__37073),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__7513 (
            .O(N__37070),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__7512 (
            .O(N__37067),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__7511 (
            .O(N__37060),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    CascadeMux I__7510 (
            .O(N__37057),
            .I(N__37054));
    InMux I__7509 (
            .O(N__37054),
            .I(N__37051));
    LocalMux I__7508 (
            .O(N__37051),
            .I(N__37047));
    InMux I__7507 (
            .O(N__37050),
            .I(N__37044));
    Span4Mux_v I__7506 (
            .O(N__37047),
            .I(N__37037));
    LocalMux I__7505 (
            .O(N__37044),
            .I(N__37037));
    InMux I__7504 (
            .O(N__37043),
            .I(N__37034));
    InMux I__7503 (
            .O(N__37042),
            .I(N__37031));
    Sp12to4 I__7502 (
            .O(N__37037),
            .I(N__37026));
    LocalMux I__7501 (
            .O(N__37034),
            .I(N__37026));
    LocalMux I__7500 (
            .O(N__37031),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv12 I__7499 (
            .O(N__37026),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__7498 (
            .O(N__37021),
            .I(N__37018));
    LocalMux I__7497 (
            .O(N__37018),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2 ));
    InMux I__7496 (
            .O(N__37015),
            .I(N__37011));
    InMux I__7495 (
            .O(N__37014),
            .I(N__37008));
    LocalMux I__7494 (
            .O(N__37011),
            .I(N__37005));
    LocalMux I__7493 (
            .O(N__37008),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__7492 (
            .O(N__37005),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__7491 (
            .O(N__37000),
            .I(N__36996));
    InMux I__7490 (
            .O(N__36999),
            .I(N__36993));
    LocalMux I__7489 (
            .O(N__36996),
            .I(N__36990));
    LocalMux I__7488 (
            .O(N__36993),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__7487 (
            .O(N__36990),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__7486 (
            .O(N__36985),
            .I(N__36982));
    LocalMux I__7485 (
            .O(N__36982),
            .I(N__36979));
    Span4Mux_h I__7484 (
            .O(N__36979),
            .I(N__36976));
    Odrv4 I__7483 (
            .O(N__36976),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df20 ));
    InMux I__7482 (
            .O(N__36973),
            .I(N__36969));
    InMux I__7481 (
            .O(N__36972),
            .I(N__36966));
    LocalMux I__7480 (
            .O(N__36969),
            .I(N__36963));
    LocalMux I__7479 (
            .O(N__36966),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__7478 (
            .O(N__36963),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__7477 (
            .O(N__36958),
            .I(N__36954));
    InMux I__7476 (
            .O(N__36957),
            .I(N__36951));
    LocalMux I__7475 (
            .O(N__36954),
            .I(N__36948));
    LocalMux I__7474 (
            .O(N__36951),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__7473 (
            .O(N__36948),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__7472 (
            .O(N__36943),
            .I(N__36940));
    LocalMux I__7471 (
            .O(N__36940),
            .I(N__36937));
    Span4Mux_h I__7470 (
            .O(N__36937),
            .I(N__36934));
    Odrv4 I__7469 (
            .O(N__36934),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df22 ));
    InMux I__7468 (
            .O(N__36931),
            .I(N__36927));
    InMux I__7467 (
            .O(N__36930),
            .I(N__36924));
    LocalMux I__7466 (
            .O(N__36927),
            .I(N__36921));
    LocalMux I__7465 (
            .O(N__36924),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__7464 (
            .O(N__36921),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__7463 (
            .O(N__36916),
            .I(N__36912));
    InMux I__7462 (
            .O(N__36915),
            .I(N__36909));
    LocalMux I__7461 (
            .O(N__36912),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    LocalMux I__7460 (
            .O(N__36909),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__7459 (
            .O(N__36904),
            .I(N__36901));
    LocalMux I__7458 (
            .O(N__36901),
            .I(N__36898));
    Span4Mux_v I__7457 (
            .O(N__36898),
            .I(N__36895));
    Odrv4 I__7456 (
            .O(N__36895),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df24 ));
    InMux I__7455 (
            .O(N__36892),
            .I(N__36888));
    InMux I__7454 (
            .O(N__36891),
            .I(N__36885));
    LocalMux I__7453 (
            .O(N__36888),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    LocalMux I__7452 (
            .O(N__36885),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    CascadeMux I__7451 (
            .O(N__36880),
            .I(N__36876));
    InMux I__7450 (
            .O(N__36879),
            .I(N__36873));
    InMux I__7449 (
            .O(N__36876),
            .I(N__36870));
    LocalMux I__7448 (
            .O(N__36873),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    LocalMux I__7447 (
            .O(N__36870),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__7446 (
            .O(N__36865),
            .I(N__36862));
    LocalMux I__7445 (
            .O(N__36862),
            .I(N__36859));
    Span4Mux_v I__7444 (
            .O(N__36859),
            .I(N__36856));
    Odrv4 I__7443 (
            .O(N__36856),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df26 ));
    InMux I__7442 (
            .O(N__36853),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__7441 (
            .O(N__36850),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__7440 (
            .O(N__36847),
            .I(bfn_14_18_0_));
    InMux I__7439 (
            .O(N__36844),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__7438 (
            .O(N__36841),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__7437 (
            .O(N__36838),
            .I(N__36835));
    LocalMux I__7436 (
            .O(N__36835),
            .I(N__36831));
    InMux I__7435 (
            .O(N__36834),
            .I(N__36828));
    Span4Mux_v I__7434 (
            .O(N__36831),
            .I(N__36825));
    LocalMux I__7433 (
            .O(N__36828),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__7432 (
            .O(N__36825),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__7431 (
            .O(N__36820),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__7430 (
            .O(N__36817),
            .I(N__36814));
    LocalMux I__7429 (
            .O(N__36814),
            .I(N__36810));
    InMux I__7428 (
            .O(N__36813),
            .I(N__36807));
    Span4Mux_v I__7427 (
            .O(N__36810),
            .I(N__36804));
    LocalMux I__7426 (
            .O(N__36807),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__7425 (
            .O(N__36804),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__7424 (
            .O(N__36799),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__7423 (
            .O(N__36796),
            .I(N__36792));
    CascadeMux I__7422 (
            .O(N__36795),
            .I(N__36789));
    LocalMux I__7421 (
            .O(N__36792),
            .I(N__36785));
    InMux I__7420 (
            .O(N__36789),
            .I(N__36782));
    InMux I__7419 (
            .O(N__36788),
            .I(N__36779));
    Span4Mux_v I__7418 (
            .O(N__36785),
            .I(N__36776));
    LocalMux I__7417 (
            .O(N__36782),
            .I(N__36773));
    LocalMux I__7416 (
            .O(N__36779),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__7415 (
            .O(N__36776),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv12 I__7414 (
            .O(N__36773),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__7413 (
            .O(N__36766),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    CEMux I__7412 (
            .O(N__36763),
            .I(N__36758));
    CEMux I__7411 (
            .O(N__36762),
            .I(N__36755));
    CEMux I__7410 (
            .O(N__36761),
            .I(N__36751));
    LocalMux I__7409 (
            .O(N__36758),
            .I(N__36740));
    LocalMux I__7408 (
            .O(N__36755),
            .I(N__36736));
    CEMux I__7407 (
            .O(N__36754),
            .I(N__36733));
    LocalMux I__7406 (
            .O(N__36751),
            .I(N__36730));
    CEMux I__7405 (
            .O(N__36750),
            .I(N__36716));
    InMux I__7404 (
            .O(N__36749),
            .I(N__36709));
    InMux I__7403 (
            .O(N__36748),
            .I(N__36709));
    InMux I__7402 (
            .O(N__36747),
            .I(N__36709));
    InMux I__7401 (
            .O(N__36746),
            .I(N__36700));
    InMux I__7400 (
            .O(N__36745),
            .I(N__36700));
    InMux I__7399 (
            .O(N__36744),
            .I(N__36700));
    InMux I__7398 (
            .O(N__36743),
            .I(N__36700));
    Span4Mux_v I__7397 (
            .O(N__36740),
            .I(N__36685));
    InMux I__7396 (
            .O(N__36739),
            .I(N__36682));
    Span4Mux_v I__7395 (
            .O(N__36736),
            .I(N__36677));
    LocalMux I__7394 (
            .O(N__36733),
            .I(N__36677));
    Span4Mux_h I__7393 (
            .O(N__36730),
            .I(N__36674));
    InMux I__7392 (
            .O(N__36729),
            .I(N__36665));
    InMux I__7391 (
            .O(N__36728),
            .I(N__36665));
    InMux I__7390 (
            .O(N__36727),
            .I(N__36665));
    InMux I__7389 (
            .O(N__36726),
            .I(N__36665));
    InMux I__7388 (
            .O(N__36725),
            .I(N__36656));
    InMux I__7387 (
            .O(N__36724),
            .I(N__36656));
    InMux I__7386 (
            .O(N__36723),
            .I(N__36656));
    InMux I__7385 (
            .O(N__36722),
            .I(N__36656));
    InMux I__7384 (
            .O(N__36721),
            .I(N__36649));
    InMux I__7383 (
            .O(N__36720),
            .I(N__36649));
    InMux I__7382 (
            .O(N__36719),
            .I(N__36649));
    LocalMux I__7381 (
            .O(N__36716),
            .I(N__36646));
    LocalMux I__7380 (
            .O(N__36709),
            .I(N__36641));
    LocalMux I__7379 (
            .O(N__36700),
            .I(N__36641));
    InMux I__7378 (
            .O(N__36699),
            .I(N__36632));
    InMux I__7377 (
            .O(N__36698),
            .I(N__36632));
    InMux I__7376 (
            .O(N__36697),
            .I(N__36632));
    InMux I__7375 (
            .O(N__36696),
            .I(N__36632));
    InMux I__7374 (
            .O(N__36695),
            .I(N__36623));
    InMux I__7373 (
            .O(N__36694),
            .I(N__36623));
    InMux I__7372 (
            .O(N__36693),
            .I(N__36623));
    InMux I__7371 (
            .O(N__36692),
            .I(N__36623));
    InMux I__7370 (
            .O(N__36691),
            .I(N__36614));
    InMux I__7369 (
            .O(N__36690),
            .I(N__36614));
    InMux I__7368 (
            .O(N__36689),
            .I(N__36614));
    InMux I__7367 (
            .O(N__36688),
            .I(N__36614));
    Span4Mux_h I__7366 (
            .O(N__36685),
            .I(N__36609));
    LocalMux I__7365 (
            .O(N__36682),
            .I(N__36609));
    Span4Mux_v I__7364 (
            .O(N__36677),
            .I(N__36606));
    Span4Mux_v I__7363 (
            .O(N__36674),
            .I(N__36601));
    LocalMux I__7362 (
            .O(N__36665),
            .I(N__36601));
    LocalMux I__7361 (
            .O(N__36656),
            .I(N__36598));
    LocalMux I__7360 (
            .O(N__36649),
            .I(N__36585));
    Span4Mux_v I__7359 (
            .O(N__36646),
            .I(N__36585));
    Span4Mux_h I__7358 (
            .O(N__36641),
            .I(N__36585));
    LocalMux I__7357 (
            .O(N__36632),
            .I(N__36585));
    LocalMux I__7356 (
            .O(N__36623),
            .I(N__36585));
    LocalMux I__7355 (
            .O(N__36614),
            .I(N__36585));
    Span4Mux_v I__7354 (
            .O(N__36609),
            .I(N__36582));
    Span4Mux_h I__7353 (
            .O(N__36606),
            .I(N__36579));
    Span4Mux_h I__7352 (
            .O(N__36601),
            .I(N__36576));
    Span4Mux_v I__7351 (
            .O(N__36598),
            .I(N__36571));
    Span4Mux_v I__7350 (
            .O(N__36585),
            .I(N__36571));
    Span4Mux_v I__7349 (
            .O(N__36582),
            .I(N__36568));
    Span4Mux_v I__7348 (
            .O(N__36579),
            .I(N__36565));
    Odrv4 I__7347 (
            .O(N__36576),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__7346 (
            .O(N__36571),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__7345 (
            .O(N__36568),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__7344 (
            .O(N__36565),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__7343 (
            .O(N__36556),
            .I(N__36552));
    InMux I__7342 (
            .O(N__36555),
            .I(N__36549));
    LocalMux I__7341 (
            .O(N__36552),
            .I(N__36546));
    LocalMux I__7340 (
            .O(N__36549),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__7339 (
            .O(N__36546),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__7338 (
            .O(N__36541),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__7337 (
            .O(N__36538),
            .I(N__36535));
    LocalMux I__7336 (
            .O(N__36535),
            .I(N__36531));
    InMux I__7335 (
            .O(N__36534),
            .I(N__36528));
    Span4Mux_v I__7334 (
            .O(N__36531),
            .I(N__36525));
    LocalMux I__7333 (
            .O(N__36528),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__7332 (
            .O(N__36525),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__7331 (
            .O(N__36520),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    CascadeMux I__7330 (
            .O(N__36517),
            .I(N__36513));
    CascadeMux I__7329 (
            .O(N__36516),
            .I(N__36510));
    InMux I__7328 (
            .O(N__36513),
            .I(N__36507));
    InMux I__7327 (
            .O(N__36510),
            .I(N__36504));
    LocalMux I__7326 (
            .O(N__36507),
            .I(N__36501));
    LocalMux I__7325 (
            .O(N__36504),
            .I(N__36497));
    Span4Mux_h I__7324 (
            .O(N__36501),
            .I(N__36494));
    InMux I__7323 (
            .O(N__36500),
            .I(N__36491));
    Span4Mux_v I__7322 (
            .O(N__36497),
            .I(N__36486));
    Span4Mux_v I__7321 (
            .O(N__36494),
            .I(N__36486));
    LocalMux I__7320 (
            .O(N__36491),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__7319 (
            .O(N__36486),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__7318 (
            .O(N__36481),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__7317 (
            .O(N__36478),
            .I(N__36474));
    InMux I__7316 (
            .O(N__36477),
            .I(N__36470));
    LocalMux I__7315 (
            .O(N__36474),
            .I(N__36467));
    InMux I__7314 (
            .O(N__36473),
            .I(N__36464));
    LocalMux I__7313 (
            .O(N__36470),
            .I(N__36461));
    Span4Mux_h I__7312 (
            .O(N__36467),
            .I(N__36458));
    LocalMux I__7311 (
            .O(N__36464),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv12 I__7310 (
            .O(N__36461),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__7309 (
            .O(N__36458),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__7308 (
            .O(N__36451),
            .I(bfn_14_17_0_));
    CascadeMux I__7307 (
            .O(N__36448),
            .I(N__36444));
    InMux I__7306 (
            .O(N__36447),
            .I(N__36439));
    InMux I__7305 (
            .O(N__36444),
            .I(N__36439));
    LocalMux I__7304 (
            .O(N__36439),
            .I(N__36435));
    InMux I__7303 (
            .O(N__36438),
            .I(N__36432));
    Span4Mux_v I__7302 (
            .O(N__36435),
            .I(N__36429));
    LocalMux I__7301 (
            .O(N__36432),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__7300 (
            .O(N__36429),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__7299 (
            .O(N__36424),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__7298 (
            .O(N__36421),
            .I(N__36414));
    InMux I__7297 (
            .O(N__36420),
            .I(N__36414));
    InMux I__7296 (
            .O(N__36419),
            .I(N__36411));
    LocalMux I__7295 (
            .O(N__36414),
            .I(N__36408));
    LocalMux I__7294 (
            .O(N__36411),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv12 I__7293 (
            .O(N__36408),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__7292 (
            .O(N__36403),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__7291 (
            .O(N__36400),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__7290 (
            .O(N__36397),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__7289 (
            .O(N__36394),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__7288 (
            .O(N__36391),
            .I(N__36388));
    LocalMux I__7287 (
            .O(N__36388),
            .I(N__36384));
    InMux I__7286 (
            .O(N__36387),
            .I(N__36381));
    Span4Mux_h I__7285 (
            .O(N__36384),
            .I(N__36378));
    LocalMux I__7284 (
            .O(N__36381),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__7283 (
            .O(N__36378),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__7282 (
            .O(N__36373),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__7281 (
            .O(N__36370),
            .I(N__36366));
    InMux I__7280 (
            .O(N__36369),
            .I(N__36363));
    LocalMux I__7279 (
            .O(N__36366),
            .I(N__36360));
    LocalMux I__7278 (
            .O(N__36363),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__7277 (
            .O(N__36360),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__7276 (
            .O(N__36355),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__7275 (
            .O(N__36352),
            .I(N__36348));
    InMux I__7274 (
            .O(N__36351),
            .I(N__36345));
    LocalMux I__7273 (
            .O(N__36348),
            .I(N__36342));
    LocalMux I__7272 (
            .O(N__36345),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__7271 (
            .O(N__36342),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__7270 (
            .O(N__36337),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__7269 (
            .O(N__36334),
            .I(N__36330));
    InMux I__7268 (
            .O(N__36333),
            .I(N__36327));
    LocalMux I__7267 (
            .O(N__36330),
            .I(N__36324));
    LocalMux I__7266 (
            .O(N__36327),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__7265 (
            .O(N__36324),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__7264 (
            .O(N__36319),
            .I(bfn_14_16_0_));
    InMux I__7263 (
            .O(N__36316),
            .I(N__36312));
    InMux I__7262 (
            .O(N__36315),
            .I(N__36309));
    LocalMux I__7261 (
            .O(N__36312),
            .I(N__36306));
    LocalMux I__7260 (
            .O(N__36309),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__7259 (
            .O(N__36306),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__7258 (
            .O(N__36301),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__7257 (
            .O(N__36298),
            .I(N__36295));
    LocalMux I__7256 (
            .O(N__36295),
            .I(N__36292));
    Span4Mux_v I__7255 (
            .O(N__36292),
            .I(N__36288));
    InMux I__7254 (
            .O(N__36291),
            .I(N__36285));
    Sp12to4 I__7253 (
            .O(N__36288),
            .I(N__36282));
    LocalMux I__7252 (
            .O(N__36285),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv12 I__7251 (
            .O(N__36282),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__7250 (
            .O(N__36277),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__7249 (
            .O(N__36274),
            .I(N__36270));
    InMux I__7248 (
            .O(N__36273),
            .I(N__36267));
    LocalMux I__7247 (
            .O(N__36270),
            .I(N__36264));
    LocalMux I__7246 (
            .O(N__36267),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__7245 (
            .O(N__36264),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__7244 (
            .O(N__36259),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__7243 (
            .O(N__36256),
            .I(N__36252));
    InMux I__7242 (
            .O(N__36255),
            .I(N__36249));
    LocalMux I__7241 (
            .O(N__36252),
            .I(N__36246));
    LocalMux I__7240 (
            .O(N__36249),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__7239 (
            .O(N__36246),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__7238 (
            .O(N__36241),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__7237 (
            .O(N__36238),
            .I(N__36235));
    LocalMux I__7236 (
            .O(N__36235),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ));
    CascadeMux I__7235 (
            .O(N__36232),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__7234 (
            .O(N__36229),
            .I(N__36225));
    InMux I__7233 (
            .O(N__36228),
            .I(N__36219));
    LocalMux I__7232 (
            .O(N__36225),
            .I(N__36216));
    InMux I__7231 (
            .O(N__36224),
            .I(N__36209));
    InMux I__7230 (
            .O(N__36223),
            .I(N__36209));
    InMux I__7229 (
            .O(N__36222),
            .I(N__36209));
    LocalMux I__7228 (
            .O(N__36219),
            .I(N__36206));
    Span4Mux_v I__7227 (
            .O(N__36216),
            .I(N__36201));
    LocalMux I__7226 (
            .O(N__36209),
            .I(N__36201));
    Span4Mux_v I__7225 (
            .O(N__36206),
            .I(N__36198));
    Span4Mux_h I__7224 (
            .O(N__36201),
            .I(N__36195));
    Odrv4 I__7223 (
            .O(N__36198),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__7222 (
            .O(N__36195),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__7221 (
            .O(N__36190),
            .I(N__36184));
    InMux I__7220 (
            .O(N__36189),
            .I(N__36184));
    LocalMux I__7219 (
            .O(N__36184),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__7218 (
            .O(N__36181),
            .I(N__36177));
    InMux I__7217 (
            .O(N__36180),
            .I(N__36174));
    LocalMux I__7216 (
            .O(N__36177),
            .I(N__36171));
    LocalMux I__7215 (
            .O(N__36174),
            .I(N__36167));
    Span4Mux_v I__7214 (
            .O(N__36171),
            .I(N__36164));
    InMux I__7213 (
            .O(N__36170),
            .I(N__36160));
    Span4Mux_h I__7212 (
            .O(N__36167),
            .I(N__36157));
    Span4Mux_h I__7211 (
            .O(N__36164),
            .I(N__36154));
    InMux I__7210 (
            .O(N__36163),
            .I(N__36151));
    LocalMux I__7209 (
            .O(N__36160),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__7208 (
            .O(N__36157),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__7207 (
            .O(N__36154),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__7206 (
            .O(N__36151),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    CascadeMux I__7205 (
            .O(N__36142),
            .I(N__36137));
    InMux I__7204 (
            .O(N__36141),
            .I(N__36132));
    InMux I__7203 (
            .O(N__36140),
            .I(N__36132));
    InMux I__7202 (
            .O(N__36137),
            .I(N__36129));
    LocalMux I__7201 (
            .O(N__36132),
            .I(N__36126));
    LocalMux I__7200 (
            .O(N__36129),
            .I(N__36122));
    Span4Mux_h I__7199 (
            .O(N__36126),
            .I(N__36119));
    InMux I__7198 (
            .O(N__36125),
            .I(N__36116));
    Odrv4 I__7197 (
            .O(N__36122),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    Odrv4 I__7196 (
            .O(N__36119),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__7195 (
            .O(N__36116),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    CascadeMux I__7194 (
            .O(N__36109),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ));
    InMux I__7193 (
            .O(N__36106),
            .I(N__36103));
    LocalMux I__7192 (
            .O(N__36103),
            .I(N__36100));
    Span4Mux_h I__7191 (
            .O(N__36100),
            .I(N__36096));
    InMux I__7190 (
            .O(N__36099),
            .I(N__36093));
    Odrv4 I__7189 (
            .O(N__36096),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__7188 (
            .O(N__36093),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    InMux I__7187 (
            .O(N__36088),
            .I(N__36085));
    LocalMux I__7186 (
            .O(N__36085),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    CascadeMux I__7185 (
            .O(N__36082),
            .I(N__36079));
    InMux I__7184 (
            .O(N__36079),
            .I(N__36075));
    CascadeMux I__7183 (
            .O(N__36078),
            .I(N__36071));
    LocalMux I__7182 (
            .O(N__36075),
            .I(N__36068));
    InMux I__7181 (
            .O(N__36074),
            .I(N__36065));
    InMux I__7180 (
            .O(N__36071),
            .I(N__36062));
    Span4Mux_h I__7179 (
            .O(N__36068),
            .I(N__36059));
    LocalMux I__7178 (
            .O(N__36065),
            .I(N__36056));
    LocalMux I__7177 (
            .O(N__36062),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__7176 (
            .O(N__36059),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__7175 (
            .O(N__36056),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__7174 (
            .O(N__36049),
            .I(N__36045));
    InMux I__7173 (
            .O(N__36048),
            .I(N__36042));
    LocalMux I__7172 (
            .O(N__36045),
            .I(N__36039));
    LocalMux I__7171 (
            .O(N__36042),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__7170 (
            .O(N__36039),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__7169 (
            .O(N__36034),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__7168 (
            .O(N__36031),
            .I(N__36028));
    InMux I__7167 (
            .O(N__36028),
            .I(N__36025));
    LocalMux I__7166 (
            .O(N__36025),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28 ));
    InMux I__7165 (
            .O(N__36022),
            .I(N__36018));
    InMux I__7164 (
            .O(N__36021),
            .I(N__36015));
    LocalMux I__7163 (
            .O(N__36018),
            .I(N__36012));
    LocalMux I__7162 (
            .O(N__36015),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__7161 (
            .O(N__36012),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__7160 (
            .O(N__36007),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__7159 (
            .O(N__36004),
            .I(N__36000));
    InMux I__7158 (
            .O(N__36003),
            .I(N__35997));
    LocalMux I__7157 (
            .O(N__36000),
            .I(N__35994));
    LocalMux I__7156 (
            .O(N__35997),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__7155 (
            .O(N__35994),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__7154 (
            .O(N__35989),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__7153 (
            .O(N__35986),
            .I(N__35982));
    InMux I__7152 (
            .O(N__35985),
            .I(N__35979));
    LocalMux I__7151 (
            .O(N__35982),
            .I(N__35976));
    LocalMux I__7150 (
            .O(N__35979),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__7149 (
            .O(N__35976),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__7148 (
            .O(N__35971),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    CascadeMux I__7147 (
            .O(N__35968),
            .I(N__35965));
    InMux I__7146 (
            .O(N__35965),
            .I(N__35962));
    LocalMux I__7145 (
            .O(N__35962),
            .I(N__35959));
    Span4Mux_v I__7144 (
            .O(N__35959),
            .I(N__35956));
    Odrv4 I__7143 (
            .O(N__35956),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    CascadeMux I__7142 (
            .O(N__35953),
            .I(N__35950));
    InMux I__7141 (
            .O(N__35950),
            .I(N__35944));
    InMux I__7140 (
            .O(N__35949),
            .I(N__35944));
    LocalMux I__7139 (
            .O(N__35944),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__7138 (
            .O(N__35941),
            .I(N__35938));
    LocalMux I__7137 (
            .O(N__35938),
            .I(N__35935));
    Odrv4 I__7136 (
            .O(N__35935),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    InMux I__7135 (
            .O(N__35932),
            .I(N__35926));
    InMux I__7134 (
            .O(N__35931),
            .I(N__35926));
    LocalMux I__7133 (
            .O(N__35926),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    InMux I__7132 (
            .O(N__35923),
            .I(N__35919));
    InMux I__7131 (
            .O(N__35922),
            .I(N__35916));
    LocalMux I__7130 (
            .O(N__35919),
            .I(N__35913));
    LocalMux I__7129 (
            .O(N__35916),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    Odrv12 I__7128 (
            .O(N__35913),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    InMux I__7127 (
            .O(N__35908),
            .I(N__35905));
    LocalMux I__7126 (
            .O(N__35905),
            .I(N__35901));
    InMux I__7125 (
            .O(N__35904),
            .I(N__35898));
    Span4Mux_v I__7124 (
            .O(N__35901),
            .I(N__35895));
    LocalMux I__7123 (
            .O(N__35898),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    Odrv4 I__7122 (
            .O(N__35895),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    InMux I__7121 (
            .O(N__35890),
            .I(N__35887));
    LocalMux I__7120 (
            .O(N__35887),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    InMux I__7119 (
            .O(N__35884),
            .I(N__35880));
    InMux I__7118 (
            .O(N__35883),
            .I(N__35877));
    LocalMux I__7117 (
            .O(N__35880),
            .I(N__35874));
    LocalMux I__7116 (
            .O(N__35877),
            .I(N__35869));
    Span12Mux_h I__7115 (
            .O(N__35874),
            .I(N__35866));
    InMux I__7114 (
            .O(N__35873),
            .I(N__35863));
    InMux I__7113 (
            .O(N__35872),
            .I(N__35860));
    Span4Mux_h I__7112 (
            .O(N__35869),
            .I(N__35857));
    Span12Mux_v I__7111 (
            .O(N__35866),
            .I(N__35854));
    LocalMux I__7110 (
            .O(N__35863),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__7109 (
            .O(N__35860),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__7108 (
            .O(N__35857),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv12 I__7107 (
            .O(N__35854),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__7106 (
            .O(N__35845),
            .I(N__35838));
    InMux I__7105 (
            .O(N__35844),
            .I(N__35838));
    InMux I__7104 (
            .O(N__35843),
            .I(N__35835));
    LocalMux I__7103 (
            .O(N__35838),
            .I(N__35832));
    LocalMux I__7102 (
            .O(N__35835),
            .I(N__35829));
    Span4Mux_v I__7101 (
            .O(N__35832),
            .I(N__35824));
    Span4Mux_h I__7100 (
            .O(N__35829),
            .I(N__35824));
    Span4Mux_h I__7099 (
            .O(N__35824),
            .I(N__35821));
    Odrv4 I__7098 (
            .O(N__35821),
            .I(il_min_comp2_D2));
    InMux I__7097 (
            .O(N__35818),
            .I(N__35814));
    InMux I__7096 (
            .O(N__35817),
            .I(N__35811));
    LocalMux I__7095 (
            .O(N__35814),
            .I(N__35808));
    LocalMux I__7094 (
            .O(N__35811),
            .I(N__35803));
    Span4Mux_v I__7093 (
            .O(N__35808),
            .I(N__35803));
    Span4Mux_v I__7092 (
            .O(N__35803),
            .I(N__35800));
    Odrv4 I__7091 (
            .O(N__35800),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    CascadeMux I__7090 (
            .O(N__35797),
            .I(\phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_ ));
    InMux I__7089 (
            .O(N__35794),
            .I(N__35790));
    InMux I__7088 (
            .O(N__35793),
            .I(N__35787));
    LocalMux I__7087 (
            .O(N__35790),
            .I(N__35784));
    LocalMux I__7086 (
            .O(N__35787),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__7085 (
            .O(N__35784),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    CascadeMux I__7084 (
            .O(N__35779),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_ ));
    InMux I__7083 (
            .O(N__35776),
            .I(N__35773));
    LocalMux I__7082 (
            .O(N__35773),
            .I(N__35769));
    InMux I__7081 (
            .O(N__35772),
            .I(N__35766));
    Odrv4 I__7080 (
            .O(N__35769),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2 ));
    LocalMux I__7079 (
            .O(N__35766),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2 ));
    CascadeMux I__7078 (
            .O(N__35761),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_ ));
    CascadeMux I__7077 (
            .O(N__35758),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_ ));
    CascadeMux I__7076 (
            .O(N__35755),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_ ));
    InMux I__7075 (
            .O(N__35752),
            .I(N__35749));
    LocalMux I__7074 (
            .O(N__35749),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    InMux I__7073 (
            .O(N__35746),
            .I(N__35743));
    LocalMux I__7072 (
            .O(N__35743),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    InMux I__7071 (
            .O(N__35740),
            .I(N__35737));
    LocalMux I__7070 (
            .O(N__35737),
            .I(N__35734));
    Span4Mux_h I__7069 (
            .O(N__35734),
            .I(N__35730));
    InMux I__7068 (
            .O(N__35733),
            .I(N__35727));
    Odrv4 I__7067 (
            .O(N__35730),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ));
    LocalMux I__7066 (
            .O(N__35727),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ));
    CascadeMux I__7065 (
            .O(N__35722),
            .I(elapsed_time_ns_1_RNIP7HF91_0_10_cascade_));
    InMux I__7064 (
            .O(N__35719),
            .I(N__35716));
    LocalMux I__7063 (
            .O(N__35716),
            .I(N__35711));
    InMux I__7062 (
            .O(N__35715),
            .I(N__35708));
    InMux I__7061 (
            .O(N__35714),
            .I(N__35704));
    Span4Mux_v I__7060 (
            .O(N__35711),
            .I(N__35701));
    LocalMux I__7059 (
            .O(N__35708),
            .I(N__35698));
    InMux I__7058 (
            .O(N__35707),
            .I(N__35695));
    LocalMux I__7057 (
            .O(N__35704),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    Odrv4 I__7056 (
            .O(N__35701),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    Odrv4 I__7055 (
            .O(N__35698),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    LocalMux I__7054 (
            .O(N__35695),
            .I(elapsed_time_ns_1_RNIFJ2591_0_7));
    CascadeMux I__7053 (
            .O(N__35686),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_ ));
    InMux I__7052 (
            .O(N__35683),
            .I(N__35680));
    LocalMux I__7051 (
            .O(N__35680),
            .I(N__35677));
    Span4Mux_v I__7050 (
            .O(N__35677),
            .I(N__35671));
    InMux I__7049 (
            .O(N__35676),
            .I(N__35668));
    InMux I__7048 (
            .O(N__35675),
            .I(N__35663));
    InMux I__7047 (
            .O(N__35674),
            .I(N__35663));
    Odrv4 I__7046 (
            .O(N__35671),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    LocalMux I__7045 (
            .O(N__35668),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    LocalMux I__7044 (
            .O(N__35663),
            .I(elapsed_time_ns_1_RNIGK2591_0_8));
    InMux I__7043 (
            .O(N__35656),
            .I(N__35652));
    InMux I__7042 (
            .O(N__35655),
            .I(N__35647));
    LocalMux I__7041 (
            .O(N__35652),
            .I(N__35644));
    InMux I__7040 (
            .O(N__35651),
            .I(N__35641));
    InMux I__7039 (
            .O(N__35650),
            .I(N__35638));
    LocalMux I__7038 (
            .O(N__35647),
            .I(N__35635));
    Span4Mux_h I__7037 (
            .O(N__35644),
            .I(N__35629));
    LocalMux I__7036 (
            .O(N__35641),
            .I(N__35629));
    LocalMux I__7035 (
            .O(N__35638),
            .I(N__35626));
    Span4Mux_v I__7034 (
            .O(N__35635),
            .I(N__35623));
    InMux I__7033 (
            .O(N__35634),
            .I(N__35620));
    Span4Mux_h I__7032 (
            .O(N__35629),
            .I(N__35617));
    Odrv12 I__7031 (
            .O(N__35626),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__7030 (
            .O(N__35623),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__7029 (
            .O(N__35620),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__7028 (
            .O(N__35617),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__7027 (
            .O(N__35608),
            .I(N__35605));
    LocalMux I__7026 (
            .O(N__35605),
            .I(N__35602));
    Odrv12 I__7025 (
            .O(N__35602),
            .I(\current_shift_inst.PI_CTRL.integrator_i_19 ));
    InMux I__7024 (
            .O(N__35599),
            .I(N__35596));
    LocalMux I__7023 (
            .O(N__35596),
            .I(N__35593));
    Span4Mux_h I__7022 (
            .O(N__35593),
            .I(N__35590));
    Odrv4 I__7021 (
            .O(N__35590),
            .I(\current_shift_inst.PI_CTRL.integrator_i_9 ));
    CascadeMux I__7020 (
            .O(N__35587),
            .I(N__35584));
    InMux I__7019 (
            .O(N__35584),
            .I(N__35580));
    InMux I__7018 (
            .O(N__35583),
            .I(N__35576));
    LocalMux I__7017 (
            .O(N__35580),
            .I(N__35573));
    InMux I__7016 (
            .O(N__35579),
            .I(N__35570));
    LocalMux I__7015 (
            .O(N__35576),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    Odrv4 I__7014 (
            .O(N__35573),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    LocalMux I__7013 (
            .O(N__35570),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ));
    CascadeMux I__7012 (
            .O(N__35563),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9_cascade_ ));
    CascadeMux I__7011 (
            .O(N__35560),
            .I(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ));
    CascadeMux I__7010 (
            .O(N__35557),
            .I(N__35554));
    InMux I__7009 (
            .O(N__35554),
            .I(N__35551));
    LocalMux I__7008 (
            .O(N__35551),
            .I(N__35548));
    Span4Mux_v I__7007 (
            .O(N__35548),
            .I(N__35545));
    Odrv4 I__7006 (
            .O(N__35545),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    InMux I__7005 (
            .O(N__35542),
            .I(N__35539));
    LocalMux I__7004 (
            .O(N__35539),
            .I(N__35536));
    Span4Mux_v I__7003 (
            .O(N__35536),
            .I(N__35533));
    Odrv4 I__7002 (
            .O(N__35533),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__7001 (
            .O(N__35530),
            .I(N__35527));
    InMux I__7000 (
            .O(N__35527),
            .I(N__35524));
    LocalMux I__6999 (
            .O(N__35524),
            .I(N__35521));
    Span4Mux_v I__6998 (
            .O(N__35521),
            .I(N__35518));
    Odrv4 I__6997 (
            .O(N__35518),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    InMux I__6996 (
            .O(N__35515),
            .I(N__35511));
    InMux I__6995 (
            .O(N__35514),
            .I(N__35507));
    LocalMux I__6994 (
            .O(N__35511),
            .I(N__35504));
    InMux I__6993 (
            .O(N__35510),
            .I(N__35501));
    LocalMux I__6992 (
            .O(N__35507),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    Odrv4 I__6991 (
            .O(N__35504),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    LocalMux I__6990 (
            .O(N__35501),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ));
    CascadeMux I__6989 (
            .O(N__35494),
            .I(N__35491));
    InMux I__6988 (
            .O(N__35491),
            .I(N__35487));
    InMux I__6987 (
            .O(N__35490),
            .I(N__35483));
    LocalMux I__6986 (
            .O(N__35487),
            .I(N__35480));
    InMux I__6985 (
            .O(N__35486),
            .I(N__35477));
    LocalMux I__6984 (
            .O(N__35483),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    Odrv4 I__6983 (
            .O(N__35480),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    LocalMux I__6982 (
            .O(N__35477),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ));
    InMux I__6981 (
            .O(N__35470),
            .I(N__35466));
    InMux I__6980 (
            .O(N__35469),
            .I(N__35463));
    LocalMux I__6979 (
            .O(N__35466),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    LocalMux I__6978 (
            .O(N__35463),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ));
    InMux I__6977 (
            .O(N__35458),
            .I(N__35453));
    InMux I__6976 (
            .O(N__35457),
            .I(N__35450));
    InMux I__6975 (
            .O(N__35456),
            .I(N__35447));
    LocalMux I__6974 (
            .O(N__35453),
            .I(N__35443));
    LocalMux I__6973 (
            .O(N__35450),
            .I(N__35439));
    LocalMux I__6972 (
            .O(N__35447),
            .I(N__35436));
    InMux I__6971 (
            .O(N__35446),
            .I(N__35433));
    Span4Mux_v I__6970 (
            .O(N__35443),
            .I(N__35430));
    InMux I__6969 (
            .O(N__35442),
            .I(N__35427));
    Span4Mux_h I__6968 (
            .O(N__35439),
            .I(N__35422));
    Span4Mux_h I__6967 (
            .O(N__35436),
            .I(N__35422));
    LocalMux I__6966 (
            .O(N__35433),
            .I(N__35419));
    Sp12to4 I__6965 (
            .O(N__35430),
            .I(N__35414));
    LocalMux I__6964 (
            .O(N__35427),
            .I(N__35414));
    Odrv4 I__6963 (
            .O(N__35422),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv12 I__6962 (
            .O(N__35419),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv12 I__6961 (
            .O(N__35414),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__6960 (
            .O(N__35407),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28_cascade_ ));
    InMux I__6959 (
            .O(N__35404),
            .I(N__35401));
    LocalMux I__6958 (
            .O(N__35401),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ));
    CascadeMux I__6957 (
            .O(N__35398),
            .I(N__35395));
    InMux I__6956 (
            .O(N__35395),
            .I(N__35392));
    LocalMux I__6955 (
            .O(N__35392),
            .I(N__35389));
    Span4Mux_h I__6954 (
            .O(N__35389),
            .I(N__35386));
    Odrv4 I__6953 (
            .O(N__35386),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0 ));
    InMux I__6952 (
            .O(N__35383),
            .I(N__35379));
    InMux I__6951 (
            .O(N__35382),
            .I(N__35376));
    LocalMux I__6950 (
            .O(N__35379),
            .I(N__35373));
    LocalMux I__6949 (
            .O(N__35376),
            .I(N__35370));
    Span4Mux_h I__6948 (
            .O(N__35373),
            .I(N__35367));
    Span4Mux_v I__6947 (
            .O(N__35370),
            .I(N__35362));
    Span4Mux_v I__6946 (
            .O(N__35367),
            .I(N__35359));
    InMux I__6945 (
            .O(N__35366),
            .I(N__35356));
    InMux I__6944 (
            .O(N__35365),
            .I(N__35353));
    Span4Mux_h I__6943 (
            .O(N__35362),
            .I(N__35348));
    Span4Mux_v I__6942 (
            .O(N__35359),
            .I(N__35348));
    LocalMux I__6941 (
            .O(N__35356),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__6940 (
            .O(N__35353),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__6939 (
            .O(N__35348),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__6938 (
            .O(N__35341),
            .I(N__35336));
    InMux I__6937 (
            .O(N__35340),
            .I(N__35333));
    InMux I__6936 (
            .O(N__35339),
            .I(N__35330));
    LocalMux I__6935 (
            .O(N__35336),
            .I(N__35327));
    LocalMux I__6934 (
            .O(N__35333),
            .I(N__35324));
    LocalMux I__6933 (
            .O(N__35330),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv4 I__6932 (
            .O(N__35327),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    Odrv4 I__6931 (
            .O(N__35324),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ));
    InMux I__6930 (
            .O(N__35317),
            .I(N__35314));
    LocalMux I__6929 (
            .O(N__35314),
            .I(N__35311));
    Odrv12 I__6928 (
            .O(N__35311),
            .I(\current_shift_inst.PI_CTRL.integrator_i_16 ));
    InMux I__6927 (
            .O(N__35308),
            .I(N__35303));
    CascadeMux I__6926 (
            .O(N__35307),
            .I(N__35300));
    InMux I__6925 (
            .O(N__35306),
            .I(N__35297));
    LocalMux I__6924 (
            .O(N__35303),
            .I(N__35294));
    InMux I__6923 (
            .O(N__35300),
            .I(N__35291));
    LocalMux I__6922 (
            .O(N__35297),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    Odrv4 I__6921 (
            .O(N__35294),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    LocalMux I__6920 (
            .O(N__35291),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ));
    CascadeMux I__6919 (
            .O(N__35284),
            .I(N__35280));
    InMux I__6918 (
            .O(N__35283),
            .I(N__35277));
    InMux I__6917 (
            .O(N__35280),
            .I(N__35274));
    LocalMux I__6916 (
            .O(N__35277),
            .I(N__35270));
    LocalMux I__6915 (
            .O(N__35274),
            .I(N__35267));
    InMux I__6914 (
            .O(N__35273),
            .I(N__35262));
    Span4Mux_v I__6913 (
            .O(N__35270),
            .I(N__35259));
    Span4Mux_v I__6912 (
            .O(N__35267),
            .I(N__35256));
    InMux I__6911 (
            .O(N__35266),
            .I(N__35251));
    InMux I__6910 (
            .O(N__35265),
            .I(N__35251));
    LocalMux I__6909 (
            .O(N__35262),
            .I(N__35248));
    Odrv4 I__6908 (
            .O(N__35259),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__6907 (
            .O(N__35256),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__6906 (
            .O(N__35251),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__6905 (
            .O(N__35248),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    CascadeMux I__6904 (
            .O(N__35239),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_ ));
    InMux I__6903 (
            .O(N__35236),
            .I(N__35233));
    LocalMux I__6902 (
            .O(N__35233),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ));
    CascadeMux I__6901 (
            .O(N__35230),
            .I(N__35227));
    InMux I__6900 (
            .O(N__35227),
            .I(N__35224));
    LocalMux I__6899 (
            .O(N__35224),
            .I(N__35221));
    Span12Mux_h I__6898 (
            .O(N__35221),
            .I(N__35218));
    Odrv12 I__6897 (
            .O(N__35218),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0 ));
    InMux I__6896 (
            .O(N__35215),
            .I(N__35212));
    LocalMux I__6895 (
            .O(N__35212),
            .I(N__35208));
    InMux I__6894 (
            .O(N__35211),
            .I(N__35204));
    Span4Mux_h I__6893 (
            .O(N__35208),
            .I(N__35201));
    InMux I__6892 (
            .O(N__35207),
            .I(N__35198));
    LocalMux I__6891 (
            .O(N__35204),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    Odrv4 I__6890 (
            .O(N__35201),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    LocalMux I__6889 (
            .O(N__35198),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ));
    CascadeMux I__6888 (
            .O(N__35191),
            .I(N__35187));
    InMux I__6887 (
            .O(N__35190),
            .I(N__35184));
    InMux I__6886 (
            .O(N__35187),
            .I(N__35180));
    LocalMux I__6885 (
            .O(N__35184),
            .I(N__35177));
    InMux I__6884 (
            .O(N__35183),
            .I(N__35174));
    LocalMux I__6883 (
            .O(N__35180),
            .I(N__35171));
    Span4Mux_h I__6882 (
            .O(N__35177),
            .I(N__35168));
    LocalMux I__6881 (
            .O(N__35174),
            .I(N__35165));
    Span4Mux_h I__6880 (
            .O(N__35171),
            .I(N__35162));
    Span4Mux_v I__6879 (
            .O(N__35168),
            .I(N__35159));
    Odrv4 I__6878 (
            .O(N__35165),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__6877 (
            .O(N__35162),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv4 I__6876 (
            .O(N__35159),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__6875 (
            .O(N__35152),
            .I(N__35149));
    LocalMux I__6874 (
            .O(N__35149),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_12 ));
    CascadeMux I__6873 (
            .O(N__35146),
            .I(N__35143));
    InMux I__6872 (
            .O(N__35143),
            .I(N__35140));
    LocalMux I__6871 (
            .O(N__35140),
            .I(N__35137));
    Span4Mux_h I__6870 (
            .O(N__35137),
            .I(N__35134));
    Odrv4 I__6869 (
            .O(N__35134),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12 ));
    InMux I__6868 (
            .O(N__35131),
            .I(N__35127));
    CascadeMux I__6867 (
            .O(N__35130),
            .I(N__35124));
    LocalMux I__6866 (
            .O(N__35127),
            .I(N__35120));
    InMux I__6865 (
            .O(N__35124),
            .I(N__35117));
    InMux I__6864 (
            .O(N__35123),
            .I(N__35114));
    Span4Mux_v I__6863 (
            .O(N__35120),
            .I(N__35111));
    LocalMux I__6862 (
            .O(N__35117),
            .I(N__35108));
    LocalMux I__6861 (
            .O(N__35114),
            .I(N__35105));
    Span4Mux_h I__6860 (
            .O(N__35111),
            .I(N__35098));
    Span4Mux_h I__6859 (
            .O(N__35108),
            .I(N__35098));
    Span4Mux_h I__6858 (
            .O(N__35105),
            .I(N__35095));
    InMux I__6857 (
            .O(N__35104),
            .I(N__35092));
    InMux I__6856 (
            .O(N__35103),
            .I(N__35089));
    Odrv4 I__6855 (
            .O(N__35098),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__6854 (
            .O(N__35095),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__6853 (
            .O(N__35092),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__6852 (
            .O(N__35089),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__6851 (
            .O(N__35080),
            .I(N__35075));
    InMux I__6850 (
            .O(N__35079),
            .I(N__35072));
    InMux I__6849 (
            .O(N__35078),
            .I(N__35069));
    LocalMux I__6848 (
            .O(N__35075),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    LocalMux I__6847 (
            .O(N__35072),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    LocalMux I__6846 (
            .O(N__35069),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ));
    InMux I__6845 (
            .O(N__35062),
            .I(N__35059));
    LocalMux I__6844 (
            .O(N__35059),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ));
    CascadeMux I__6843 (
            .O(N__35056),
            .I(N__35053));
    InMux I__6842 (
            .O(N__35053),
            .I(N__35050));
    LocalMux I__6841 (
            .O(N__35050),
            .I(N__35047));
    Span4Mux_h I__6840 (
            .O(N__35047),
            .I(N__35044));
    Odrv4 I__6839 (
            .O(N__35044),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0 ));
    InMux I__6838 (
            .O(N__35041),
            .I(N__35037));
    InMux I__6837 (
            .O(N__35040),
            .I(N__35033));
    LocalMux I__6836 (
            .O(N__35037),
            .I(N__35030));
    InMux I__6835 (
            .O(N__35036),
            .I(N__35027));
    LocalMux I__6834 (
            .O(N__35033),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    Odrv4 I__6833 (
            .O(N__35030),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    LocalMux I__6832 (
            .O(N__35027),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ));
    InMux I__6831 (
            .O(N__35020),
            .I(N__35015));
    InMux I__6830 (
            .O(N__35019),
            .I(N__35012));
    InMux I__6829 (
            .O(N__35018),
            .I(N__35009));
    LocalMux I__6828 (
            .O(N__35015),
            .I(N__35004));
    LocalMux I__6827 (
            .O(N__35012),
            .I(N__35004));
    LocalMux I__6826 (
            .O(N__35009),
            .I(N__35001));
    Span4Mux_h I__6825 (
            .O(N__35004),
            .I(N__34998));
    Odrv12 I__6824 (
            .O(N__35001),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__6823 (
            .O(N__34998),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__6822 (
            .O(N__34993),
            .I(N__34990));
    LocalMux I__6821 (
            .O(N__34990),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ));
    InMux I__6820 (
            .O(N__34987),
            .I(N__34984));
    LocalMux I__6819 (
            .O(N__34984),
            .I(N__34980));
    InMux I__6818 (
            .O(N__34983),
            .I(N__34976));
    Span4Mux_h I__6817 (
            .O(N__34980),
            .I(N__34973));
    InMux I__6816 (
            .O(N__34979),
            .I(N__34970));
    LocalMux I__6815 (
            .O(N__34976),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    Odrv4 I__6814 (
            .O(N__34973),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    LocalMux I__6813 (
            .O(N__34970),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ));
    CascadeMux I__6812 (
            .O(N__34963),
            .I(N__34958));
    InMux I__6811 (
            .O(N__34962),
            .I(N__34950));
    InMux I__6810 (
            .O(N__34961),
            .I(N__34950));
    InMux I__6809 (
            .O(N__34958),
            .I(N__34950));
    InMux I__6808 (
            .O(N__34957),
            .I(N__34947));
    LocalMux I__6807 (
            .O(N__34950),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__6806 (
            .O(N__34947),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    IoInMux I__6805 (
            .O(N__34942),
            .I(N__34939));
    LocalMux I__6804 (
            .O(N__34939),
            .I(N__34936));
    Span12Mux_s6_v I__6803 (
            .O(N__34936),
            .I(N__34931));
    InMux I__6802 (
            .O(N__34935),
            .I(N__34926));
    InMux I__6801 (
            .O(N__34934),
            .I(N__34926));
    Odrv12 I__6800 (
            .O(N__34931),
            .I(s1_phy_c));
    LocalMux I__6799 (
            .O(N__34926),
            .I(s1_phy_c));
    InMux I__6798 (
            .O(N__34921),
            .I(N__34915));
    InMux I__6797 (
            .O(N__34920),
            .I(N__34910));
    InMux I__6796 (
            .O(N__34919),
            .I(N__34910));
    InMux I__6795 (
            .O(N__34918),
            .I(N__34907));
    LocalMux I__6794 (
            .O(N__34915),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__6793 (
            .O(N__34910),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__6792 (
            .O(N__34907),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    IoInMux I__6791 (
            .O(N__34900),
            .I(N__34897));
    LocalMux I__6790 (
            .O(N__34897),
            .I(N__34894));
    Span4Mux_s3_v I__6789 (
            .O(N__34894),
            .I(N__34891));
    Span4Mux_h I__6788 (
            .O(N__34891),
            .I(N__34887));
    InMux I__6787 (
            .O(N__34890),
            .I(N__34884));
    Odrv4 I__6786 (
            .O(N__34887),
            .I(T23_c));
    LocalMux I__6785 (
            .O(N__34884),
            .I(T23_c));
    InMux I__6784 (
            .O(N__34879),
            .I(N__34874));
    InMux I__6783 (
            .O(N__34878),
            .I(N__34870));
    InMux I__6782 (
            .O(N__34877),
            .I(N__34867));
    LocalMux I__6781 (
            .O(N__34874),
            .I(N__34864));
    InMux I__6780 (
            .O(N__34873),
            .I(N__34861));
    LocalMux I__6779 (
            .O(N__34870),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__6778 (
            .O(N__34867),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv12 I__6777 (
            .O(N__34864),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__6776 (
            .O(N__34861),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__6775 (
            .O(N__34852),
            .I(N__34844));
    InMux I__6774 (
            .O(N__34851),
            .I(N__34844));
    InMux I__6773 (
            .O(N__34850),
            .I(N__34841));
    InMux I__6772 (
            .O(N__34849),
            .I(N__34838));
    LocalMux I__6771 (
            .O(N__34844),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6770 (
            .O(N__34841),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__6769 (
            .O(N__34838),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__6768 (
            .O(N__34831),
            .I(N__34828));
    LocalMux I__6767 (
            .O(N__34828),
            .I(N__34825));
    Odrv12 I__6766 (
            .O(N__34825),
            .I(\current_shift_inst.timer_s1.N_166_i ));
    IoInMux I__6765 (
            .O(N__34822),
            .I(N__34819));
    LocalMux I__6764 (
            .O(N__34819),
            .I(N__34816));
    Odrv12 I__6763 (
            .O(N__34816),
            .I(s2_phy_c));
    InMux I__6762 (
            .O(N__34813),
            .I(N__34810));
    LocalMux I__6761 (
            .O(N__34810),
            .I(N__34807));
    Span4Mux_h I__6760 (
            .O(N__34807),
            .I(N__34804));
    Odrv4 I__6759 (
            .O(N__34804),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    CascadeMux I__6758 (
            .O(N__34801),
            .I(N__34798));
    InMux I__6757 (
            .O(N__34798),
            .I(N__34793));
    InMux I__6756 (
            .O(N__34797),
            .I(N__34790));
    InMux I__6755 (
            .O(N__34796),
            .I(N__34787));
    LocalMux I__6754 (
            .O(N__34793),
            .I(N__34784));
    LocalMux I__6753 (
            .O(N__34790),
            .I(N__34779));
    LocalMux I__6752 (
            .O(N__34787),
            .I(N__34779));
    Span4Mux_v I__6751 (
            .O(N__34784),
            .I(N__34776));
    Span4Mux_v I__6750 (
            .O(N__34779),
            .I(N__34771));
    Span4Mux_v I__6749 (
            .O(N__34776),
            .I(N__34768));
    InMux I__6748 (
            .O(N__34775),
            .I(N__34763));
    InMux I__6747 (
            .O(N__34774),
            .I(N__34763));
    Sp12to4 I__6746 (
            .O(N__34771),
            .I(N__34756));
    Sp12to4 I__6745 (
            .O(N__34768),
            .I(N__34756));
    LocalMux I__6744 (
            .O(N__34763),
            .I(N__34756));
    Odrv12 I__6743 (
            .O(N__34756),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__6742 (
            .O(N__34753),
            .I(N__34750));
    LocalMux I__6741 (
            .O(N__34750),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ));
    InMux I__6740 (
            .O(N__34747),
            .I(N__34743));
    InMux I__6739 (
            .O(N__34746),
            .I(N__34740));
    LocalMux I__6738 (
            .O(N__34743),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    LocalMux I__6737 (
            .O(N__34740),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ));
    InMux I__6736 (
            .O(N__34735),
            .I(N__34731));
    InMux I__6735 (
            .O(N__34734),
            .I(N__34728));
    LocalMux I__6734 (
            .O(N__34731),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ));
    LocalMux I__6733 (
            .O(N__34728),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ));
    CascadeMux I__6732 (
            .O(N__34723),
            .I(elapsed_time_ns_1_RNIP93CP1_0_1_cascade_));
    CascadeMux I__6731 (
            .O(N__34720),
            .I(N__34716));
    InMux I__6730 (
            .O(N__34719),
            .I(N__34713));
    InMux I__6729 (
            .O(N__34716),
            .I(N__34710));
    LocalMux I__6728 (
            .O(N__34713),
            .I(N__34705));
    LocalMux I__6727 (
            .O(N__34710),
            .I(N__34705));
    Odrv4 I__6726 (
            .O(N__34705),
            .I(\phase_controller_inst1.stoper_hc.N_310 ));
    CascadeMux I__6725 (
            .O(N__34702),
            .I(N__34698));
    InMux I__6724 (
            .O(N__34701),
            .I(N__34695));
    InMux I__6723 (
            .O(N__34698),
            .I(N__34692));
    LocalMux I__6722 (
            .O(N__34695),
            .I(N__34689));
    LocalMux I__6721 (
            .O(N__34692),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ));
    Odrv4 I__6720 (
            .O(N__34689),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ));
    CascadeMux I__6719 (
            .O(N__34684),
            .I(N__34681));
    InMux I__6718 (
            .O(N__34681),
            .I(N__34678));
    LocalMux I__6717 (
            .O(N__34678),
            .I(N__34675));
    Odrv4 I__6716 (
            .O(N__34675),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__6715 (
            .O(N__34672),
            .I(N__34668));
    InMux I__6714 (
            .O(N__34671),
            .I(N__34665));
    LocalMux I__6713 (
            .O(N__34668),
            .I(state_ns_i_a2_1));
    LocalMux I__6712 (
            .O(N__34665),
            .I(state_ns_i_a2_1));
    InMux I__6711 (
            .O(N__34660),
            .I(N__34656));
    InMux I__6710 (
            .O(N__34659),
            .I(N__34653));
    LocalMux I__6709 (
            .O(N__34656),
            .I(N__34650));
    LocalMux I__6708 (
            .O(N__34653),
            .I(N__34646));
    Span4Mux_v I__6707 (
            .O(N__34650),
            .I(N__34643));
    InMux I__6706 (
            .O(N__34649),
            .I(N__34640));
    Span12Mux_s9_v I__6705 (
            .O(N__34646),
            .I(N__34637));
    Odrv4 I__6704 (
            .O(N__34643),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__6703 (
            .O(N__34640),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv12 I__6702 (
            .O(N__34637),
            .I(\phase_controller_inst1.tr_time_passed ));
    IoInMux I__6701 (
            .O(N__34630),
            .I(N__34627));
    LocalMux I__6700 (
            .O(N__34627),
            .I(N__34624));
    Span4Mux_s3_v I__6699 (
            .O(N__34624),
            .I(N__34621));
    Span4Mux_v I__6698 (
            .O(N__34621),
            .I(N__34617));
    InMux I__6697 (
            .O(N__34620),
            .I(N__34614));
    Odrv4 I__6696 (
            .O(N__34617),
            .I(T45_c));
    LocalMux I__6695 (
            .O(N__34614),
            .I(T45_c));
    CascadeMux I__6694 (
            .O(N__34609),
            .I(N__34604));
    InMux I__6693 (
            .O(N__34608),
            .I(N__34601));
    CascadeMux I__6692 (
            .O(N__34607),
            .I(N__34598));
    InMux I__6691 (
            .O(N__34604),
            .I(N__34594));
    LocalMux I__6690 (
            .O(N__34601),
            .I(N__34591));
    InMux I__6689 (
            .O(N__34598),
            .I(N__34588));
    InMux I__6688 (
            .O(N__34597),
            .I(N__34585));
    LocalMux I__6687 (
            .O(N__34594),
            .I(elapsed_time_ns_1_RNIRB3CP1_0_3));
    Odrv4 I__6686 (
            .O(N__34591),
            .I(elapsed_time_ns_1_RNIRB3CP1_0_3));
    LocalMux I__6685 (
            .O(N__34588),
            .I(elapsed_time_ns_1_RNIRB3CP1_0_3));
    LocalMux I__6684 (
            .O(N__34585),
            .I(elapsed_time_ns_1_RNIRB3CP1_0_3));
    CascadeMux I__6683 (
            .O(N__34576),
            .I(N__34573));
    InMux I__6682 (
            .O(N__34573),
            .I(N__34564));
    InMux I__6681 (
            .O(N__34572),
            .I(N__34564));
    InMux I__6680 (
            .O(N__34571),
            .I(N__34564));
    LocalMux I__6679 (
            .O(N__34564),
            .I(elapsed_time_ns_1_RNIJEKEE1_0_2));
    InMux I__6678 (
            .O(N__34561),
            .I(N__34558));
    LocalMux I__6677 (
            .O(N__34558),
            .I(\phase_controller_inst1.stoper_hc.N_286 ));
    CascadeMux I__6676 (
            .O(N__34555),
            .I(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1_cascade_ ));
    InMux I__6675 (
            .O(N__34552),
            .I(N__34546));
    InMux I__6674 (
            .O(N__34551),
            .I(N__34546));
    LocalMux I__6673 (
            .O(N__34546),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    CascadeMux I__6672 (
            .O(N__34543),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_ ));
    CascadeMux I__6671 (
            .O(N__34540),
            .I(\phase_controller_inst1.stoper_hc.N_328_cascade_ ));
    CascadeMux I__6670 (
            .O(N__34537),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ));
    InMux I__6669 (
            .O(N__34534),
            .I(N__34529));
    InMux I__6668 (
            .O(N__34533),
            .I(N__34524));
    InMux I__6667 (
            .O(N__34532),
            .I(N__34524));
    LocalMux I__6666 (
            .O(N__34529),
            .I(elapsed_time_ns_1_RNIP93CP1_0_1));
    LocalMux I__6665 (
            .O(N__34524),
            .I(elapsed_time_ns_1_RNIP93CP1_0_1));
    InMux I__6664 (
            .O(N__34519),
            .I(N__34515));
    InMux I__6663 (
            .O(N__34518),
            .I(N__34512));
    LocalMux I__6662 (
            .O(N__34515),
            .I(N__34507));
    LocalMux I__6661 (
            .O(N__34512),
            .I(N__34507));
    Span4Mux_v I__6660 (
            .O(N__34507),
            .I(N__34502));
    InMux I__6659 (
            .O(N__34506),
            .I(N__34497));
    InMux I__6658 (
            .O(N__34505),
            .I(N__34497));
    Odrv4 I__6657 (
            .O(N__34502),
            .I(elapsed_time_ns_1_RNIPKKEE1_0_8));
    LocalMux I__6656 (
            .O(N__34497),
            .I(elapsed_time_ns_1_RNIPKKEE1_0_8));
    CascadeMux I__6655 (
            .O(N__34492),
            .I(elapsed_time_ns_1_RNIOJKEE1_0_7_cascade_));
    CascadeMux I__6654 (
            .O(N__34489),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ));
    CascadeMux I__6653 (
            .O(N__34486),
            .I(\phase_controller_inst1.stoper_hc.N_330_cascade_ ));
    InMux I__6652 (
            .O(N__34483),
            .I(N__34479));
    InMux I__6651 (
            .O(N__34482),
            .I(N__34476));
    LocalMux I__6650 (
            .O(N__34479),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ));
    LocalMux I__6649 (
            .O(N__34476),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ));
    InMux I__6648 (
            .O(N__34471),
            .I(N__34467));
    InMux I__6647 (
            .O(N__34470),
            .I(N__34464));
    LocalMux I__6646 (
            .O(N__34467),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2 ));
    LocalMux I__6645 (
            .O(N__34464),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2 ));
    CascadeMux I__6644 (
            .O(N__34459),
            .I(N__34456));
    InMux I__6643 (
            .O(N__34456),
            .I(N__34451));
    InMux I__6642 (
            .O(N__34455),
            .I(N__34446));
    InMux I__6641 (
            .O(N__34454),
            .I(N__34446));
    LocalMux I__6640 (
            .O(N__34451),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ));
    LocalMux I__6639 (
            .O(N__34446),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ));
    CascadeMux I__6638 (
            .O(N__34441),
            .I(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_ ));
    InMux I__6637 (
            .O(N__34438),
            .I(N__34435));
    LocalMux I__6636 (
            .O(N__34435),
            .I(N__34432));
    Odrv12 I__6635 (
            .O(N__34432),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df28 ));
    InMux I__6634 (
            .O(N__34429),
            .I(N__34426));
    LocalMux I__6633 (
            .O(N__34426),
            .I(N__34423));
    Odrv12 I__6632 (
            .O(N__34423),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    InMux I__6631 (
            .O(N__34420),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ));
    InMux I__6630 (
            .O(N__34417),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    CascadeMux I__6629 (
            .O(N__34414),
            .I(N__34411));
    InMux I__6628 (
            .O(N__34411),
            .I(N__34408));
    LocalMux I__6627 (
            .O(N__34408),
            .I(N__34405));
    Odrv12 I__6626 (
            .O(N__34405),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    InMux I__6625 (
            .O(N__34402),
            .I(N__34399));
    LocalMux I__6624 (
            .O(N__34399),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__6623 (
            .O(N__34396),
            .I(N__34393));
    LocalMux I__6622 (
            .O(N__34393),
            .I(N__34390));
    Odrv12 I__6621 (
            .O(N__34390),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__6620 (
            .O(N__34387),
            .I(N__34384));
    InMux I__6619 (
            .O(N__34384),
            .I(N__34381));
    LocalMux I__6618 (
            .O(N__34381),
            .I(N__34378));
    Odrv4 I__6617 (
            .O(N__34378),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__6616 (
            .O(N__34375),
            .I(N__34372));
    LocalMux I__6615 (
            .O(N__34372),
            .I(N__34369));
    Odrv12 I__6614 (
            .O(N__34369),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__6613 (
            .O(N__34366),
            .I(N__34363));
    InMux I__6612 (
            .O(N__34363),
            .I(N__34360));
    LocalMux I__6611 (
            .O(N__34360),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__6610 (
            .O(N__34357),
            .I(N__34354));
    LocalMux I__6609 (
            .O(N__34354),
            .I(N__34351));
    Odrv12 I__6608 (
            .O(N__34351),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__6607 (
            .O(N__34348),
            .I(N__34345));
    InMux I__6606 (
            .O(N__34345),
            .I(N__34342));
    LocalMux I__6605 (
            .O(N__34342),
            .I(N__34339));
    Odrv4 I__6604 (
            .O(N__34339),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__6603 (
            .O(N__34336),
            .I(N__34333));
    LocalMux I__6602 (
            .O(N__34333),
            .I(N__34330));
    Odrv12 I__6601 (
            .O(N__34330),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__6600 (
            .O(N__34327),
            .I(N__34324));
    InMux I__6599 (
            .O(N__34324),
            .I(N__34321));
    LocalMux I__6598 (
            .O(N__34321),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__6597 (
            .O(N__34318),
            .I(N__34315));
    InMux I__6596 (
            .O(N__34315),
            .I(N__34312));
    LocalMux I__6595 (
            .O(N__34312),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    CascadeMux I__6594 (
            .O(N__34309),
            .I(N__34306));
    InMux I__6593 (
            .O(N__34306),
            .I(N__34303));
    LocalMux I__6592 (
            .O(N__34303),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__6591 (
            .O(N__34300),
            .I(N__34297));
    LocalMux I__6590 (
            .O(N__34297),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__6589 (
            .O(N__34294),
            .I(N__34291));
    InMux I__6588 (
            .O(N__34291),
            .I(N__34288));
    LocalMux I__6587 (
            .O(N__34288),
            .I(N__34285));
    Odrv4 I__6586 (
            .O(N__34285),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__6585 (
            .O(N__34282),
            .I(N__34279));
    LocalMux I__6584 (
            .O(N__34279),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__6583 (
            .O(N__34276),
            .I(N__34273));
    InMux I__6582 (
            .O(N__34273),
            .I(N__34270));
    LocalMux I__6581 (
            .O(N__34270),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__6580 (
            .O(N__34267),
            .I(N__34264));
    LocalMux I__6579 (
            .O(N__34264),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__6578 (
            .O(N__34261),
            .I(N__34258));
    InMux I__6577 (
            .O(N__34258),
            .I(N__34255));
    LocalMux I__6576 (
            .O(N__34255),
            .I(N__34252));
    Odrv4 I__6575 (
            .O(N__34252),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__6574 (
            .O(N__34249),
            .I(N__34246));
    LocalMux I__6573 (
            .O(N__34246),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__6572 (
            .O(N__34243),
            .I(N__34240));
    InMux I__6571 (
            .O(N__34240),
            .I(N__34237));
    LocalMux I__6570 (
            .O(N__34237),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__6569 (
            .O(N__34234),
            .I(N__34231));
    InMux I__6568 (
            .O(N__34231),
            .I(N__34228));
    LocalMux I__6567 (
            .O(N__34228),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    InMux I__6566 (
            .O(N__34225),
            .I(N__34222));
    LocalMux I__6565 (
            .O(N__34222),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    CascadeMux I__6564 (
            .O(N__34219),
            .I(N__34216));
    InMux I__6563 (
            .O(N__34216),
            .I(N__34213));
    LocalMux I__6562 (
            .O(N__34213),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    InMux I__6561 (
            .O(N__34210),
            .I(N__34207));
    LocalMux I__6560 (
            .O(N__34207),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__6559 (
            .O(N__34204),
            .I(N__34201));
    LocalMux I__6558 (
            .O(N__34201),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    IoInMux I__6557 (
            .O(N__34198),
            .I(N__34195));
    LocalMux I__6556 (
            .O(N__34195),
            .I(N__34192));
    IoSpan4Mux I__6555 (
            .O(N__34192),
            .I(N__34189));
    Span4Mux_s1_v I__6554 (
            .O(N__34189),
            .I(N__34186));
    Sp12to4 I__6553 (
            .O(N__34186),
            .I(N__34183));
    Span12Mux_s9_v I__6552 (
            .O(N__34183),
            .I(N__34180));
    Odrv12 I__6551 (
            .O(N__34180),
            .I(\pll_inst.red_c_i ));
    InMux I__6550 (
            .O(N__34177),
            .I(N__34174));
    LocalMux I__6549 (
            .O(N__34174),
            .I(N__34169));
    InMux I__6548 (
            .O(N__34173),
            .I(N__34166));
    InMux I__6547 (
            .O(N__34172),
            .I(N__34163));
    Sp12to4 I__6546 (
            .O(N__34169),
            .I(N__34158));
    LocalMux I__6545 (
            .O(N__34166),
            .I(N__34158));
    LocalMux I__6544 (
            .O(N__34163),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    Odrv12 I__6543 (
            .O(N__34158),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ));
    CascadeMux I__6542 (
            .O(N__34153),
            .I(N__34150));
    InMux I__6541 (
            .O(N__34150),
            .I(N__34147));
    LocalMux I__6540 (
            .O(N__34147),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__6539 (
            .O(N__34144),
            .I(N__34141));
    LocalMux I__6538 (
            .O(N__34141),
            .I(N__34136));
    InMux I__6537 (
            .O(N__34140),
            .I(N__34133));
    InMux I__6536 (
            .O(N__34139),
            .I(N__34130));
    Sp12to4 I__6535 (
            .O(N__34136),
            .I(N__34125));
    LocalMux I__6534 (
            .O(N__34133),
            .I(N__34125));
    LocalMux I__6533 (
            .O(N__34130),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    Odrv12 I__6532 (
            .O(N__34125),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ));
    InMux I__6531 (
            .O(N__34120),
            .I(N__34117));
    LocalMux I__6530 (
            .O(N__34117),
            .I(N__34114));
    Odrv4 I__6529 (
            .O(N__34114),
            .I(\current_shift_inst.PI_CTRL.integrator_i_24 ));
    InMux I__6528 (
            .O(N__34111),
            .I(N__34106));
    InMux I__6527 (
            .O(N__34110),
            .I(N__34103));
    InMux I__6526 (
            .O(N__34109),
            .I(N__34100));
    LocalMux I__6525 (
            .O(N__34106),
            .I(N__34097));
    LocalMux I__6524 (
            .O(N__34103),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    LocalMux I__6523 (
            .O(N__34100),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    Odrv12 I__6522 (
            .O(N__34097),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ));
    CascadeMux I__6521 (
            .O(N__34090),
            .I(N__34087));
    InMux I__6520 (
            .O(N__34087),
            .I(N__34081));
    InMux I__6519 (
            .O(N__34086),
            .I(N__34078));
    InMux I__6518 (
            .O(N__34085),
            .I(N__34075));
    InMux I__6517 (
            .O(N__34084),
            .I(N__34072));
    LocalMux I__6516 (
            .O(N__34081),
            .I(N__34069));
    LocalMux I__6515 (
            .O(N__34078),
            .I(N__34066));
    LocalMux I__6514 (
            .O(N__34075),
            .I(N__34061));
    LocalMux I__6513 (
            .O(N__34072),
            .I(N__34061));
    Span4Mux_h I__6512 (
            .O(N__34069),
            .I(N__34057));
    Span4Mux_v I__6511 (
            .O(N__34066),
            .I(N__34052));
    Span4Mux_v I__6510 (
            .O(N__34061),
            .I(N__34052));
    InMux I__6509 (
            .O(N__34060),
            .I(N__34049));
    Odrv4 I__6508 (
            .O(N__34057),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__6507 (
            .O(N__34052),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__6506 (
            .O(N__34049),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__6505 (
            .O(N__34042),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_31 ));
    InMux I__6504 (
            .O(N__34039),
            .I(N__34036));
    LocalMux I__6503 (
            .O(N__34036),
            .I(N__34033));
    Span4Mux_h I__6502 (
            .O(N__34033),
            .I(N__34030));
    Odrv4 I__6501 (
            .O(N__34030),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0 ));
    CascadeMux I__6500 (
            .O(N__34027),
            .I(N__34024));
    InMux I__6499 (
            .O(N__34024),
            .I(N__34021));
    LocalMux I__6498 (
            .O(N__34021),
            .I(N__34018));
    Odrv12 I__6497 (
            .O(N__34018),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    CascadeMux I__6496 (
            .O(N__34015),
            .I(N__34012));
    InMux I__6495 (
            .O(N__34012),
            .I(N__34008));
    CascadeMux I__6494 (
            .O(N__34011),
            .I(N__34003));
    LocalMux I__6493 (
            .O(N__34008),
            .I(N__33999));
    InMux I__6492 (
            .O(N__34007),
            .I(N__33994));
    InMux I__6491 (
            .O(N__34006),
            .I(N__33994));
    InMux I__6490 (
            .O(N__34003),
            .I(N__33989));
    InMux I__6489 (
            .O(N__34002),
            .I(N__33989));
    Span12Mux_v I__6488 (
            .O(N__33999),
            .I(N__33984));
    LocalMux I__6487 (
            .O(N__33994),
            .I(N__33984));
    LocalMux I__6486 (
            .O(N__33989),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv12 I__6485 (
            .O(N__33984),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__6484 (
            .O(N__33979),
            .I(N__33976));
    InMux I__6483 (
            .O(N__33976),
            .I(N__33973));
    LocalMux I__6482 (
            .O(N__33973),
            .I(N__33970));
    Odrv4 I__6481 (
            .O(N__33970),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__6480 (
            .O(N__33967),
            .I(N__33964));
    LocalMux I__6479 (
            .O(N__33964),
            .I(N__33961));
    Span4Mux_h I__6478 (
            .O(N__33961),
            .I(N__33958));
    Odrv4 I__6477 (
            .O(N__33958),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    CascadeMux I__6476 (
            .O(N__33955),
            .I(N__33952));
    InMux I__6475 (
            .O(N__33952),
            .I(N__33946));
    InMux I__6474 (
            .O(N__33951),
            .I(N__33943));
    InMux I__6473 (
            .O(N__33950),
            .I(N__33940));
    InMux I__6472 (
            .O(N__33949),
            .I(N__33937));
    LocalMux I__6471 (
            .O(N__33946),
            .I(N__33933));
    LocalMux I__6470 (
            .O(N__33943),
            .I(N__33930));
    LocalMux I__6469 (
            .O(N__33940),
            .I(N__33927));
    LocalMux I__6468 (
            .O(N__33937),
            .I(N__33924));
    InMux I__6467 (
            .O(N__33936),
            .I(N__33921));
    Span4Mux_v I__6466 (
            .O(N__33933),
            .I(N__33918));
    Span4Mux_v I__6465 (
            .O(N__33930),
            .I(N__33911));
    Span4Mux_v I__6464 (
            .O(N__33927),
            .I(N__33911));
    Span4Mux_v I__6463 (
            .O(N__33924),
            .I(N__33911));
    LocalMux I__6462 (
            .O(N__33921),
            .I(N__33908));
    Span4Mux_h I__6461 (
            .O(N__33918),
            .I(N__33905));
    Span4Mux_h I__6460 (
            .O(N__33911),
            .I(N__33902));
    Odrv12 I__6459 (
            .O(N__33908),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__6458 (
            .O(N__33905),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__6457 (
            .O(N__33902),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    CascadeMux I__6456 (
            .O(N__33895),
            .I(N__33892));
    InMux I__6455 (
            .O(N__33892),
            .I(N__33889));
    LocalMux I__6454 (
            .O(N__33889),
            .I(N__33886));
    Odrv4 I__6453 (
            .O(N__33886),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__6452 (
            .O(N__33883),
            .I(N__33880));
    LocalMux I__6451 (
            .O(N__33880),
            .I(N__33877));
    Span4Mux_h I__6450 (
            .O(N__33877),
            .I(N__33874));
    Odrv4 I__6449 (
            .O(N__33874),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__6448 (
            .O(N__33871),
            .I(N__33868));
    InMux I__6447 (
            .O(N__33868),
            .I(N__33864));
    InMux I__6446 (
            .O(N__33867),
            .I(N__33859));
    LocalMux I__6445 (
            .O(N__33864),
            .I(N__33856));
    InMux I__6444 (
            .O(N__33863),
            .I(N__33853));
    InMux I__6443 (
            .O(N__33862),
            .I(N__33850));
    LocalMux I__6442 (
            .O(N__33859),
            .I(N__33847));
    Span4Mux_v I__6441 (
            .O(N__33856),
            .I(N__33844));
    LocalMux I__6440 (
            .O(N__33853),
            .I(N__33841));
    LocalMux I__6439 (
            .O(N__33850),
            .I(N__33837));
    Span4Mux_v I__6438 (
            .O(N__33847),
            .I(N__33832));
    Span4Mux_h I__6437 (
            .O(N__33844),
            .I(N__33832));
    Span4Mux_v I__6436 (
            .O(N__33841),
            .I(N__33829));
    InMux I__6435 (
            .O(N__33840),
            .I(N__33826));
    Odrv12 I__6434 (
            .O(N__33837),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__6433 (
            .O(N__33832),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__6432 (
            .O(N__33829),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__6431 (
            .O(N__33826),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    InMux I__6430 (
            .O(N__33817),
            .I(N__33814));
    LocalMux I__6429 (
            .O(N__33814),
            .I(N__33809));
    CascadeMux I__6428 (
            .O(N__33813),
            .I(N__33806));
    CascadeMux I__6427 (
            .O(N__33812),
            .I(N__33803));
    Span4Mux_h I__6426 (
            .O(N__33809),
            .I(N__33799));
    InMux I__6425 (
            .O(N__33806),
            .I(N__33796));
    InMux I__6424 (
            .O(N__33803),
            .I(N__33793));
    InMux I__6423 (
            .O(N__33802),
            .I(N__33789));
    Span4Mux_h I__6422 (
            .O(N__33799),
            .I(N__33786));
    LocalMux I__6421 (
            .O(N__33796),
            .I(N__33781));
    LocalMux I__6420 (
            .O(N__33793),
            .I(N__33781));
    InMux I__6419 (
            .O(N__33792),
            .I(N__33778));
    LocalMux I__6418 (
            .O(N__33789),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__6417 (
            .O(N__33786),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv12 I__6416 (
            .O(N__33781),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__6415 (
            .O(N__33778),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    CascadeMux I__6414 (
            .O(N__33769),
            .I(N__33766));
    InMux I__6413 (
            .O(N__33766),
            .I(N__33763));
    LocalMux I__6412 (
            .O(N__33763),
            .I(N__33760));
    Span4Mux_v I__6411 (
            .O(N__33760),
            .I(N__33757));
    Odrv4 I__6410 (
            .O(N__33757),
            .I(\current_shift_inst.PI_CTRL.integrator_i_21 ));
    CascadeMux I__6409 (
            .O(N__33754),
            .I(N__33750));
    InMux I__6408 (
            .O(N__33753),
            .I(N__33747));
    InMux I__6407 (
            .O(N__33750),
            .I(N__33744));
    LocalMux I__6406 (
            .O(N__33747),
            .I(N__33740));
    LocalMux I__6405 (
            .O(N__33744),
            .I(N__33737));
    InMux I__6404 (
            .O(N__33743),
            .I(N__33734));
    Odrv4 I__6403 (
            .O(N__33740),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv12 I__6402 (
            .O(N__33737),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    LocalMux I__6401 (
            .O(N__33734),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__6400 (
            .O(N__33727),
            .I(N__33724));
    LocalMux I__6399 (
            .O(N__33724),
            .I(N__33721));
    Odrv12 I__6398 (
            .O(N__33721),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ));
    InMux I__6397 (
            .O(N__33718),
            .I(N__33713));
    InMux I__6396 (
            .O(N__33717),
            .I(N__33710));
    InMux I__6395 (
            .O(N__33716),
            .I(N__33707));
    LocalMux I__6394 (
            .O(N__33713),
            .I(N__33704));
    LocalMux I__6393 (
            .O(N__33710),
            .I(N__33699));
    LocalMux I__6392 (
            .O(N__33707),
            .I(N__33696));
    Span4Mux_h I__6391 (
            .O(N__33704),
            .I(N__33693));
    InMux I__6390 (
            .O(N__33703),
            .I(N__33688));
    InMux I__6389 (
            .O(N__33702),
            .I(N__33688));
    Span4Mux_h I__6388 (
            .O(N__33699),
            .I(N__33685));
    Odrv4 I__6387 (
            .O(N__33696),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__6386 (
            .O(N__33693),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__6385 (
            .O(N__33688),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__6384 (
            .O(N__33685),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__6383 (
            .O(N__33676),
            .I(N__33673));
    LocalMux I__6382 (
            .O(N__33673),
            .I(N__33670));
    Span4Mux_h I__6381 (
            .O(N__33670),
            .I(N__33667));
    Odrv4 I__6380 (
            .O(N__33667),
            .I(\current_shift_inst.PI_CTRL.integrator_i_17 ));
    CascadeMux I__6379 (
            .O(N__33664),
            .I(N__33661));
    InMux I__6378 (
            .O(N__33661),
            .I(N__33658));
    LocalMux I__6377 (
            .O(N__33658),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ));
    InMux I__6376 (
            .O(N__33655),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ));
    InMux I__6375 (
            .O(N__33652),
            .I(N__33649));
    LocalMux I__6374 (
            .O(N__33649),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ));
    InMux I__6373 (
            .O(N__33646),
            .I(bfn_13_7_0_));
    InMux I__6372 (
            .O(N__33643),
            .I(N__33639));
    InMux I__6371 (
            .O(N__33642),
            .I(N__33636));
    LocalMux I__6370 (
            .O(N__33639),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    LocalMux I__6369 (
            .O(N__33636),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ));
    InMux I__6368 (
            .O(N__33631),
            .I(N__33628));
    LocalMux I__6367 (
            .O(N__33628),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ));
    InMux I__6366 (
            .O(N__33625),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ));
    InMux I__6365 (
            .O(N__33622),
            .I(N__33619));
    LocalMux I__6364 (
            .O(N__33619),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ));
    InMux I__6363 (
            .O(N__33616),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ));
    InMux I__6362 (
            .O(N__33613),
            .I(N__33610));
    LocalMux I__6361 (
            .O(N__33610),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ));
    InMux I__6360 (
            .O(N__33607),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ));
    InMux I__6359 (
            .O(N__33604),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ));
    InMux I__6358 (
            .O(N__33601),
            .I(N__33598));
    LocalMux I__6357 (
            .O(N__33598),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ));
    InMux I__6356 (
            .O(N__33595),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ));
    InMux I__6355 (
            .O(N__33592),
            .I(N__33589));
    LocalMux I__6354 (
            .O(N__33589),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ));
    InMux I__6353 (
            .O(N__33586),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ));
    CascadeMux I__6352 (
            .O(N__33583),
            .I(N__33580));
    InMux I__6351 (
            .O(N__33580),
            .I(N__33577));
    LocalMux I__6350 (
            .O(N__33577),
            .I(N__33574));
    Odrv4 I__6349 (
            .O(N__33574),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ));
    InMux I__6348 (
            .O(N__33571),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ));
    InMux I__6347 (
            .O(N__33568),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ));
    InMux I__6346 (
            .O(N__33565),
            .I(N__33562));
    LocalMux I__6345 (
            .O(N__33562),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ));
    InMux I__6344 (
            .O(N__33559),
            .I(bfn_13_6_0_));
    InMux I__6343 (
            .O(N__33556),
            .I(N__33553));
    LocalMux I__6342 (
            .O(N__33553),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ));
    InMux I__6341 (
            .O(N__33550),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ));
    InMux I__6340 (
            .O(N__33547),
            .I(N__33542));
    InMux I__6339 (
            .O(N__33546),
            .I(N__33539));
    InMux I__6338 (
            .O(N__33545),
            .I(N__33536));
    LocalMux I__6337 (
            .O(N__33542),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    LocalMux I__6336 (
            .O(N__33539),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    LocalMux I__6335 (
            .O(N__33536),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ));
    CascadeMux I__6334 (
            .O(N__33529),
            .I(N__33526));
    InMux I__6333 (
            .O(N__33526),
            .I(N__33523));
    LocalMux I__6332 (
            .O(N__33523),
            .I(N__33520));
    Odrv4 I__6331 (
            .O(N__33520),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ));
    InMux I__6330 (
            .O(N__33517),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ));
    CascadeMux I__6329 (
            .O(N__33514),
            .I(N__33511));
    InMux I__6328 (
            .O(N__33511),
            .I(N__33508));
    LocalMux I__6327 (
            .O(N__33508),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ));
    InMux I__6326 (
            .O(N__33505),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ));
    InMux I__6325 (
            .O(N__33502),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ));
    InMux I__6324 (
            .O(N__33499),
            .I(N__33496));
    LocalMux I__6323 (
            .O(N__33496),
            .I(N__33493));
    Odrv4 I__6322 (
            .O(N__33493),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ));
    InMux I__6321 (
            .O(N__33490),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ));
    InMux I__6320 (
            .O(N__33487),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ));
    InMux I__6319 (
            .O(N__33484),
            .I(N__33481));
    LocalMux I__6318 (
            .O(N__33481),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ));
    InMux I__6317 (
            .O(N__33478),
            .I(N__33475));
    LocalMux I__6316 (
            .O(N__33475),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_6 ));
    InMux I__6315 (
            .O(N__33472),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ));
    InMux I__6314 (
            .O(N__33469),
            .I(N__33466));
    LocalMux I__6313 (
            .O(N__33466),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ));
    CascadeMux I__6312 (
            .O(N__33463),
            .I(N__33460));
    InMux I__6311 (
            .O(N__33460),
            .I(N__33457));
    LocalMux I__6310 (
            .O(N__33457),
            .I(N__33454));
    Odrv4 I__6309 (
            .O(N__33454),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_7 ));
    InMux I__6308 (
            .O(N__33451),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ));
    InMux I__6307 (
            .O(N__33448),
            .I(N__33445));
    LocalMux I__6306 (
            .O(N__33445),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ));
    InMux I__6305 (
            .O(N__33442),
            .I(N__33439));
    LocalMux I__6304 (
            .O(N__33439),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_8 ));
    InMux I__6303 (
            .O(N__33436),
            .I(bfn_13_5_0_));
    CascadeMux I__6302 (
            .O(N__33433),
            .I(N__33430));
    InMux I__6301 (
            .O(N__33430),
            .I(N__33427));
    LocalMux I__6300 (
            .O(N__33427),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_9 ));
    InMux I__6299 (
            .O(N__33424),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ));
    InMux I__6298 (
            .O(N__33421),
            .I(N__33418));
    LocalMux I__6297 (
            .O(N__33418),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ));
    CascadeMux I__6296 (
            .O(N__33415),
            .I(N__33412));
    InMux I__6295 (
            .O(N__33412),
            .I(N__33409));
    LocalMux I__6294 (
            .O(N__33409),
            .I(N__33406));
    Odrv4 I__6293 (
            .O(N__33406),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_10 ));
    InMux I__6292 (
            .O(N__33403),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ));
    InMux I__6291 (
            .O(N__33400),
            .I(N__33397));
    LocalMux I__6290 (
            .O(N__33397),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ));
    CascadeMux I__6289 (
            .O(N__33394),
            .I(N__33391));
    InMux I__6288 (
            .O(N__33391),
            .I(N__33388));
    LocalMux I__6287 (
            .O(N__33388),
            .I(N__33385));
    Odrv4 I__6286 (
            .O(N__33385),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_11 ));
    InMux I__6285 (
            .O(N__33382),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ));
    InMux I__6284 (
            .O(N__33379),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ));
    InMux I__6283 (
            .O(N__33376),
            .I(N__33373));
    LocalMux I__6282 (
            .O(N__33373),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_13 ));
    InMux I__6281 (
            .O(N__33370),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ));
    InMux I__6280 (
            .O(N__33367),
            .I(N__33361));
    InMux I__6279 (
            .O(N__33366),
            .I(N__33361));
    LocalMux I__6278 (
            .O(N__33361),
            .I(\phase_controller_inst1.N_54 ));
    CEMux I__6277 (
            .O(N__33358),
            .I(N__33353));
    CEMux I__6276 (
            .O(N__33357),
            .I(N__33350));
    CEMux I__6275 (
            .O(N__33356),
            .I(N__33347));
    LocalMux I__6274 (
            .O(N__33353),
            .I(N__33342));
    LocalMux I__6273 (
            .O(N__33350),
            .I(N__33342));
    LocalMux I__6272 (
            .O(N__33347),
            .I(N__33338));
    Span4Mux_v I__6271 (
            .O(N__33342),
            .I(N__33335));
    CEMux I__6270 (
            .O(N__33341),
            .I(N__33332));
    Span4Mux_v I__6269 (
            .O(N__33338),
            .I(N__33325));
    Span4Mux_h I__6268 (
            .O(N__33335),
            .I(N__33325));
    LocalMux I__6267 (
            .O(N__33332),
            .I(N__33325));
    Span4Mux_h I__6266 (
            .O(N__33325),
            .I(N__33322));
    Span4Mux_h I__6265 (
            .O(N__33322),
            .I(N__33319));
    Odrv4 I__6264 (
            .O(N__33319),
            .I(\current_shift_inst.timer_s1.N_167_i ));
    InMux I__6263 (
            .O(N__33316),
            .I(N__33313));
    LocalMux I__6262 (
            .O(N__33313),
            .I(N__33309));
    InMux I__6261 (
            .O(N__33312),
            .I(N__33306));
    Span4Mux_h I__6260 (
            .O(N__33309),
            .I(N__33303));
    LocalMux I__6259 (
            .O(N__33306),
            .I(N__33298));
    Span4Mux_v I__6258 (
            .O(N__33303),
            .I(N__33298));
    Odrv4 I__6257 (
            .O(N__33298),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__6256 (
            .O(N__33295),
            .I(N__33292));
    LocalMux I__6255 (
            .O(N__33292),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ));
    InMux I__6254 (
            .O(N__33289),
            .I(N__33285));
    InMux I__6253 (
            .O(N__33288),
            .I(N__33282));
    LocalMux I__6252 (
            .O(N__33285),
            .I(N__33279));
    LocalMux I__6251 (
            .O(N__33282),
            .I(N__33276));
    Span4Mux_v I__6250 (
            .O(N__33279),
            .I(N__33273));
    Odrv4 I__6249 (
            .O(N__33276),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    Odrv4 I__6248 (
            .O(N__33273),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    CascadeMux I__6247 (
            .O(N__33268),
            .I(N__33265));
    InMux I__6246 (
            .O(N__33265),
            .I(N__33262));
    LocalMux I__6245 (
            .O(N__33262),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ));
    InMux I__6244 (
            .O(N__33259),
            .I(N__33255));
    InMux I__6243 (
            .O(N__33258),
            .I(N__33252));
    LocalMux I__6242 (
            .O(N__33255),
            .I(N__33249));
    LocalMux I__6241 (
            .O(N__33252),
            .I(N__33246));
    Span4Mux_v I__6240 (
            .O(N__33249),
            .I(N__33243));
    Odrv4 I__6239 (
            .O(N__33246),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv4 I__6238 (
            .O(N__33243),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__6237 (
            .O(N__33238),
            .I(N__33235));
    LocalMux I__6236 (
            .O(N__33235),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ));
    InMux I__6235 (
            .O(N__33232),
            .I(N__33228));
    InMux I__6234 (
            .O(N__33231),
            .I(N__33225));
    LocalMux I__6233 (
            .O(N__33228),
            .I(N__33222));
    LocalMux I__6232 (
            .O(N__33225),
            .I(N__33219));
    Span4Mux_v I__6231 (
            .O(N__33222),
            .I(N__33216));
    Odrv12 I__6230 (
            .O(N__33219),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv4 I__6229 (
            .O(N__33216),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__6228 (
            .O(N__33211),
            .I(N__33208));
    LocalMux I__6227 (
            .O(N__33208),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ));
    InMux I__6226 (
            .O(N__33205),
            .I(N__33202));
    LocalMux I__6225 (
            .O(N__33202),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ));
    InMux I__6224 (
            .O(N__33199),
            .I(N__33196));
    LocalMux I__6223 (
            .O(N__33196),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_4 ));
    InMux I__6222 (
            .O(N__33193),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ));
    InMux I__6221 (
            .O(N__33190),
            .I(N__33187));
    LocalMux I__6220 (
            .O(N__33187),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ));
    InMux I__6219 (
            .O(N__33184),
            .I(N__33181));
    LocalMux I__6218 (
            .O(N__33181),
            .I(\current_shift_inst.PI_CTRL.un7_integrator1_5 ));
    InMux I__6217 (
            .O(N__33178),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ));
    CascadeMux I__6216 (
            .O(N__33175),
            .I(N__33172));
    InMux I__6215 (
            .O(N__33172),
            .I(N__33169));
    LocalMux I__6214 (
            .O(N__33169),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__6213 (
            .O(N__33166),
            .I(N__33163));
    LocalMux I__6212 (
            .O(N__33163),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__6211 (
            .O(N__33160),
            .I(N__33157));
    LocalMux I__6210 (
            .O(N__33157),
            .I(N__33153));
    InMux I__6209 (
            .O(N__33156),
            .I(N__33150));
    Span4Mux_s1_v I__6208 (
            .O(N__33153),
            .I(N__33144));
    LocalMux I__6207 (
            .O(N__33150),
            .I(N__33144));
    InMux I__6206 (
            .O(N__33149),
            .I(N__33141));
    Span4Mux_v I__6205 (
            .O(N__33144),
            .I(N__33137));
    LocalMux I__6204 (
            .O(N__33141),
            .I(N__33134));
    InMux I__6203 (
            .O(N__33140),
            .I(N__33131));
    Span4Mux_h I__6202 (
            .O(N__33137),
            .I(N__33128));
    Span4Mux_v I__6201 (
            .O(N__33134),
            .I(N__33123));
    LocalMux I__6200 (
            .O(N__33131),
            .I(N__33123));
    Sp12to4 I__6199 (
            .O(N__33128),
            .I(N__33120));
    Span4Mux_v I__6198 (
            .O(N__33123),
            .I(N__33117));
    Span12Mux_v I__6197 (
            .O(N__33120),
            .I(N__33114));
    Span4Mux_v I__6196 (
            .O(N__33117),
            .I(N__33111));
    Span12Mux_v I__6195 (
            .O(N__33114),
            .I(N__33108));
    Sp12to4 I__6194 (
            .O(N__33111),
            .I(N__33105));
    Span12Mux_h I__6193 (
            .O(N__33108),
            .I(N__33102));
    Span12Mux_h I__6192 (
            .O(N__33105),
            .I(N__33099));
    Odrv12 I__6191 (
            .O(N__33102),
            .I(start_stop_c));
    Odrv12 I__6190 (
            .O(N__33099),
            .I(start_stop_c));
    InMux I__6189 (
            .O(N__33094),
            .I(N__33091));
    LocalMux I__6188 (
            .O(N__33091),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    InMux I__6187 (
            .O(N__33088),
            .I(N__33081));
    InMux I__6186 (
            .O(N__33087),
            .I(N__33072));
    InMux I__6185 (
            .O(N__33086),
            .I(N__33072));
    InMux I__6184 (
            .O(N__33085),
            .I(N__33072));
    InMux I__6183 (
            .O(N__33084),
            .I(N__33072));
    LocalMux I__6182 (
            .O(N__33081),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__6181 (
            .O(N__33072),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    CascadeMux I__6180 (
            .O(N__33067),
            .I(N__33063));
    InMux I__6179 (
            .O(N__33066),
            .I(N__33056));
    InMux I__6178 (
            .O(N__33063),
            .I(N__33056));
    InMux I__6177 (
            .O(N__33062),
            .I(N__33053));
    InMux I__6176 (
            .O(N__33061),
            .I(N__33050));
    LocalMux I__6175 (
            .O(N__33056),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__6174 (
            .O(N__33053),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__6173 (
            .O(N__33050),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__6172 (
            .O(N__33043),
            .I(N__33040));
    LocalMux I__6171 (
            .O(N__33040),
            .I(N__33037));
    Span4Mux_v I__6170 (
            .O(N__33037),
            .I(N__33034));
    Odrv4 I__6169 (
            .O(N__33034),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__6168 (
            .O(N__33031),
            .I(N__33028));
    LocalMux I__6167 (
            .O(N__33028),
            .I(N__33025));
    Odrv4 I__6166 (
            .O(N__33025),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__6165 (
            .O(N__33022),
            .I(N__33019));
    LocalMux I__6164 (
            .O(N__33019),
            .I(N__33016));
    Sp12to4 I__6163 (
            .O(N__33016),
            .I(N__33013));
    Odrv12 I__6162 (
            .O(N__33013),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__6161 (
            .O(N__33010),
            .I(N__33007));
    LocalMux I__6160 (
            .O(N__33007),
            .I(N__33004));
    Span4Mux_v I__6159 (
            .O(N__33004),
            .I(N__33001));
    Odrv4 I__6158 (
            .O(N__33001),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__6157 (
            .O(N__32998),
            .I(N__32995));
    LocalMux I__6156 (
            .O(N__32995),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__6155 (
            .O(N__32992),
            .I(N__32989));
    LocalMux I__6154 (
            .O(N__32989),
            .I(N__32986));
    Odrv12 I__6153 (
            .O(N__32986),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__6152 (
            .O(N__32983),
            .I(N__32980));
    LocalMux I__6151 (
            .O(N__32980),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    CascadeMux I__6150 (
            .O(N__32977),
            .I(N__32974));
    InMux I__6149 (
            .O(N__32974),
            .I(N__32971));
    LocalMux I__6148 (
            .O(N__32971),
            .I(N__32968));
    Span4Mux_v I__6147 (
            .O(N__32968),
            .I(N__32965));
    Odrv4 I__6146 (
            .O(N__32965),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__6145 (
            .O(N__32962),
            .I(N__32959));
    LocalMux I__6144 (
            .O(N__32959),
            .I(N__32956));
    Odrv12 I__6143 (
            .O(N__32956),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__6142 (
            .O(N__32953),
            .I(N__32950));
    LocalMux I__6141 (
            .O(N__32950),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__6140 (
            .O(N__32947),
            .I(N__32944));
    LocalMux I__6139 (
            .O(N__32944),
            .I(N__32941));
    Span4Mux_h I__6138 (
            .O(N__32941),
            .I(N__32938));
    Odrv4 I__6137 (
            .O(N__32938),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__6136 (
            .O(N__32935),
            .I(N__32932));
    LocalMux I__6135 (
            .O(N__32932),
            .I(N__32929));
    Span12Mux_h I__6134 (
            .O(N__32929),
            .I(N__32926));
    Odrv12 I__6133 (
            .O(N__32926),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__6132 (
            .O(N__32923),
            .I(N__32920));
    LocalMux I__6131 (
            .O(N__32920),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__6130 (
            .O(N__32917),
            .I(N__32914));
    LocalMux I__6129 (
            .O(N__32914),
            .I(N__32911));
    Span4Mux_h I__6128 (
            .O(N__32911),
            .I(N__32908));
    Odrv4 I__6127 (
            .O(N__32908),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__6126 (
            .O(N__32905),
            .I(N__32902));
    LocalMux I__6125 (
            .O(N__32902),
            .I(N__32899));
    Span12Mux_s11_v I__6124 (
            .O(N__32899),
            .I(N__32896));
    Odrv12 I__6123 (
            .O(N__32896),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__6122 (
            .O(N__32893),
            .I(N__32888));
    InMux I__6121 (
            .O(N__32892),
            .I(N__32885));
    InMux I__6120 (
            .O(N__32891),
            .I(N__32882));
    LocalMux I__6119 (
            .O(N__32888),
            .I(N__32878));
    LocalMux I__6118 (
            .O(N__32885),
            .I(N__32873));
    LocalMux I__6117 (
            .O(N__32882),
            .I(N__32873));
    InMux I__6116 (
            .O(N__32881),
            .I(N__32870));
    Span12Mux_v I__6115 (
            .O(N__32878),
            .I(N__32867));
    Span12Mux_v I__6114 (
            .O(N__32873),
            .I(N__32864));
    LocalMux I__6113 (
            .O(N__32870),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__6112 (
            .O(N__32867),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__6111 (
            .O(N__32864),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__6110 (
            .O(N__32857),
            .I(N__32854));
    LocalMux I__6109 (
            .O(N__32854),
            .I(N__32845));
    InMux I__6108 (
            .O(N__32853),
            .I(N__32842));
    InMux I__6107 (
            .O(N__32852),
            .I(N__32835));
    InMux I__6106 (
            .O(N__32851),
            .I(N__32835));
    InMux I__6105 (
            .O(N__32850),
            .I(N__32835));
    CascadeMux I__6104 (
            .O(N__32849),
            .I(N__32832));
    InMux I__6103 (
            .O(N__32848),
            .I(N__32829));
    Span4Mux_h I__6102 (
            .O(N__32845),
            .I(N__32814));
    LocalMux I__6101 (
            .O(N__32842),
            .I(N__32814));
    LocalMux I__6100 (
            .O(N__32835),
            .I(N__32814));
    InMux I__6099 (
            .O(N__32832),
            .I(N__32811));
    LocalMux I__6098 (
            .O(N__32829),
            .I(N__32808));
    InMux I__6097 (
            .O(N__32828),
            .I(N__32805));
    InMux I__6096 (
            .O(N__32827),
            .I(N__32790));
    InMux I__6095 (
            .O(N__32826),
            .I(N__32790));
    InMux I__6094 (
            .O(N__32825),
            .I(N__32790));
    InMux I__6093 (
            .O(N__32824),
            .I(N__32790));
    InMux I__6092 (
            .O(N__32823),
            .I(N__32790));
    InMux I__6091 (
            .O(N__32822),
            .I(N__32790));
    InMux I__6090 (
            .O(N__32821),
            .I(N__32790));
    Span4Mux_h I__6089 (
            .O(N__32814),
            .I(N__32787));
    LocalMux I__6088 (
            .O(N__32811),
            .I(N__32778));
    Span4Mux_v I__6087 (
            .O(N__32808),
            .I(N__32778));
    LocalMux I__6086 (
            .O(N__32805),
            .I(N__32778));
    LocalMux I__6085 (
            .O(N__32790),
            .I(N__32778));
    Span4Mux_v I__6084 (
            .O(N__32787),
            .I(N__32775));
    Span4Mux_v I__6083 (
            .O(N__32778),
            .I(N__32770));
    Span4Mux_v I__6082 (
            .O(N__32775),
            .I(N__32770));
    Odrv4 I__6081 (
            .O(N__32770),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__6080 (
            .O(N__32767),
            .I(N__32764));
    LocalMux I__6079 (
            .O(N__32764),
            .I(N__32761));
    Span4Mux_h I__6078 (
            .O(N__32761),
            .I(N__32758));
    Odrv4 I__6077 (
            .O(N__32758),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__6076 (
            .O(N__32755),
            .I(N__32752));
    LocalMux I__6075 (
            .O(N__32752),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__6074 (
            .O(N__32749),
            .I(N__32746));
    LocalMux I__6073 (
            .O(N__32746),
            .I(N__32743));
    Span4Mux_h I__6072 (
            .O(N__32743),
            .I(N__32740));
    Span4Mux_v I__6071 (
            .O(N__32740),
            .I(N__32737));
    Odrv4 I__6070 (
            .O(N__32737),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__6069 (
            .O(N__32734),
            .I(N__32731));
    LocalMux I__6068 (
            .O(N__32731),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__6067 (
            .O(N__32728),
            .I(N__32712));
    CascadeMux I__6066 (
            .O(N__32727),
            .I(N__32708));
    CascadeMux I__6065 (
            .O(N__32726),
            .I(N__32705));
    CascadeMux I__6064 (
            .O(N__32725),
            .I(N__32702));
    CascadeMux I__6063 (
            .O(N__32724),
            .I(N__32697));
    CascadeMux I__6062 (
            .O(N__32723),
            .I(N__32694));
    InMux I__6061 (
            .O(N__32722),
            .I(N__32678));
    InMux I__6060 (
            .O(N__32721),
            .I(N__32678));
    InMux I__6059 (
            .O(N__32720),
            .I(N__32678));
    InMux I__6058 (
            .O(N__32719),
            .I(N__32678));
    InMux I__6057 (
            .O(N__32718),
            .I(N__32678));
    InMux I__6056 (
            .O(N__32717),
            .I(N__32678));
    InMux I__6055 (
            .O(N__32716),
            .I(N__32678));
    CascadeMux I__6054 (
            .O(N__32715),
            .I(N__32674));
    InMux I__6053 (
            .O(N__32712),
            .I(N__32662));
    InMux I__6052 (
            .O(N__32711),
            .I(N__32662));
    InMux I__6051 (
            .O(N__32708),
            .I(N__32655));
    InMux I__6050 (
            .O(N__32705),
            .I(N__32655));
    InMux I__6049 (
            .O(N__32702),
            .I(N__32655));
    InMux I__6048 (
            .O(N__32701),
            .I(N__32622));
    InMux I__6047 (
            .O(N__32700),
            .I(N__32622));
    InMux I__6046 (
            .O(N__32697),
            .I(N__32622));
    InMux I__6045 (
            .O(N__32694),
            .I(N__32622));
    InMux I__6044 (
            .O(N__32693),
            .I(N__32622));
    LocalMux I__6043 (
            .O(N__32678),
            .I(N__32619));
    InMux I__6042 (
            .O(N__32677),
            .I(N__32610));
    InMux I__6041 (
            .O(N__32674),
            .I(N__32610));
    InMux I__6040 (
            .O(N__32673),
            .I(N__32610));
    InMux I__6039 (
            .O(N__32672),
            .I(N__32610));
    CascadeMux I__6038 (
            .O(N__32671),
            .I(N__32607));
    CascadeMux I__6037 (
            .O(N__32670),
            .I(N__32603));
    CascadeMux I__6036 (
            .O(N__32669),
            .I(N__32599));
    CascadeMux I__6035 (
            .O(N__32668),
            .I(N__32589));
    InMux I__6034 (
            .O(N__32667),
            .I(N__32582));
    LocalMux I__6033 (
            .O(N__32662),
            .I(N__32579));
    LocalMux I__6032 (
            .O(N__32655),
            .I(N__32576));
    CascadeMux I__6031 (
            .O(N__32654),
            .I(N__32573));
    CascadeMux I__6030 (
            .O(N__32653),
            .I(N__32566));
    CascadeMux I__6029 (
            .O(N__32652),
            .I(N__32562));
    CascadeMux I__6028 (
            .O(N__32651),
            .I(N__32558));
    CascadeMux I__6027 (
            .O(N__32650),
            .I(N__32554));
    CascadeMux I__6026 (
            .O(N__32649),
            .I(N__32550));
    CascadeMux I__6025 (
            .O(N__32648),
            .I(N__32546));
    CascadeMux I__6024 (
            .O(N__32647),
            .I(N__32542));
    CascadeMux I__6023 (
            .O(N__32646),
            .I(N__32538));
    InMux I__6022 (
            .O(N__32645),
            .I(N__32507));
    InMux I__6021 (
            .O(N__32644),
            .I(N__32507));
    InMux I__6020 (
            .O(N__32643),
            .I(N__32507));
    InMux I__6019 (
            .O(N__32642),
            .I(N__32507));
    InMux I__6018 (
            .O(N__32641),
            .I(N__32507));
    InMux I__6017 (
            .O(N__32640),
            .I(N__32507));
    InMux I__6016 (
            .O(N__32639),
            .I(N__32507));
    InMux I__6015 (
            .O(N__32638),
            .I(N__32494));
    InMux I__6014 (
            .O(N__32637),
            .I(N__32494));
    InMux I__6013 (
            .O(N__32636),
            .I(N__32494));
    InMux I__6012 (
            .O(N__32635),
            .I(N__32494));
    InMux I__6011 (
            .O(N__32634),
            .I(N__32494));
    InMux I__6010 (
            .O(N__32633),
            .I(N__32494));
    LocalMux I__6009 (
            .O(N__32622),
            .I(N__32487));
    Span4Mux_v I__6008 (
            .O(N__32619),
            .I(N__32487));
    LocalMux I__6007 (
            .O(N__32610),
            .I(N__32487));
    InMux I__6006 (
            .O(N__32607),
            .I(N__32474));
    InMux I__6005 (
            .O(N__32606),
            .I(N__32474));
    InMux I__6004 (
            .O(N__32603),
            .I(N__32474));
    InMux I__6003 (
            .O(N__32602),
            .I(N__32474));
    InMux I__6002 (
            .O(N__32599),
            .I(N__32474));
    InMux I__6001 (
            .O(N__32598),
            .I(N__32474));
    InMux I__6000 (
            .O(N__32597),
            .I(N__32461));
    InMux I__5999 (
            .O(N__32596),
            .I(N__32461));
    InMux I__5998 (
            .O(N__32595),
            .I(N__32461));
    InMux I__5997 (
            .O(N__32594),
            .I(N__32461));
    InMux I__5996 (
            .O(N__32593),
            .I(N__32461));
    InMux I__5995 (
            .O(N__32592),
            .I(N__32461));
    InMux I__5994 (
            .O(N__32589),
            .I(N__32458));
    CascadeMux I__5993 (
            .O(N__32588),
            .I(N__32448));
    CascadeMux I__5992 (
            .O(N__32587),
            .I(N__32440));
    CascadeMux I__5991 (
            .O(N__32586),
            .I(N__32436));
    CascadeMux I__5990 (
            .O(N__32585),
            .I(N__32432));
    LocalMux I__5989 (
            .O(N__32582),
            .I(N__32428));
    Span4Mux_v I__5988 (
            .O(N__32579),
            .I(N__32423));
    Span4Mux_v I__5987 (
            .O(N__32576),
            .I(N__32423));
    InMux I__5986 (
            .O(N__32573),
            .I(N__32410));
    InMux I__5985 (
            .O(N__32572),
            .I(N__32410));
    InMux I__5984 (
            .O(N__32571),
            .I(N__32410));
    InMux I__5983 (
            .O(N__32570),
            .I(N__32410));
    InMux I__5982 (
            .O(N__32569),
            .I(N__32410));
    InMux I__5981 (
            .O(N__32566),
            .I(N__32410));
    InMux I__5980 (
            .O(N__32565),
            .I(N__32395));
    InMux I__5979 (
            .O(N__32562),
            .I(N__32395));
    InMux I__5978 (
            .O(N__32561),
            .I(N__32395));
    InMux I__5977 (
            .O(N__32558),
            .I(N__32395));
    InMux I__5976 (
            .O(N__32557),
            .I(N__32395));
    InMux I__5975 (
            .O(N__32554),
            .I(N__32395));
    InMux I__5974 (
            .O(N__32553),
            .I(N__32395));
    InMux I__5973 (
            .O(N__32550),
            .I(N__32378));
    InMux I__5972 (
            .O(N__32549),
            .I(N__32378));
    InMux I__5971 (
            .O(N__32546),
            .I(N__32378));
    InMux I__5970 (
            .O(N__32545),
            .I(N__32378));
    InMux I__5969 (
            .O(N__32542),
            .I(N__32378));
    InMux I__5968 (
            .O(N__32541),
            .I(N__32378));
    InMux I__5967 (
            .O(N__32538),
            .I(N__32378));
    InMux I__5966 (
            .O(N__32537),
            .I(N__32378));
    CascadeMux I__5965 (
            .O(N__32536),
            .I(N__32375));
    CascadeMux I__5964 (
            .O(N__32535),
            .I(N__32371));
    CascadeMux I__5963 (
            .O(N__32534),
            .I(N__32367));
    CascadeMux I__5962 (
            .O(N__32533),
            .I(N__32363));
    CascadeMux I__5961 (
            .O(N__32532),
            .I(N__32359));
    CascadeMux I__5960 (
            .O(N__32531),
            .I(N__32355));
    CascadeMux I__5959 (
            .O(N__32530),
            .I(N__32351));
    CascadeMux I__5958 (
            .O(N__32529),
            .I(N__32347));
    CascadeMux I__5957 (
            .O(N__32528),
            .I(N__32343));
    CascadeMux I__5956 (
            .O(N__32527),
            .I(N__32339));
    CascadeMux I__5955 (
            .O(N__32526),
            .I(N__32335));
    CascadeMux I__5954 (
            .O(N__32525),
            .I(N__32331));
    CascadeMux I__5953 (
            .O(N__32524),
            .I(N__32327));
    CascadeMux I__5952 (
            .O(N__32523),
            .I(N__32323));
    CascadeMux I__5951 (
            .O(N__32522),
            .I(N__32319));
    LocalMux I__5950 (
            .O(N__32507),
            .I(N__32309));
    LocalMux I__5949 (
            .O(N__32494),
            .I(N__32309));
    Span4Mux_v I__5948 (
            .O(N__32487),
            .I(N__32309));
    LocalMux I__5947 (
            .O(N__32474),
            .I(N__32309));
    LocalMux I__5946 (
            .O(N__32461),
            .I(N__32306));
    LocalMux I__5945 (
            .O(N__32458),
            .I(N__32303));
    InMux I__5944 (
            .O(N__32457),
            .I(N__32288));
    InMux I__5943 (
            .O(N__32456),
            .I(N__32288));
    InMux I__5942 (
            .O(N__32455),
            .I(N__32288));
    InMux I__5941 (
            .O(N__32454),
            .I(N__32288));
    InMux I__5940 (
            .O(N__32453),
            .I(N__32288));
    InMux I__5939 (
            .O(N__32452),
            .I(N__32288));
    InMux I__5938 (
            .O(N__32451),
            .I(N__32288));
    InMux I__5937 (
            .O(N__32448),
            .I(N__32281));
    InMux I__5936 (
            .O(N__32447),
            .I(N__32281));
    InMux I__5935 (
            .O(N__32446),
            .I(N__32281));
    InMux I__5934 (
            .O(N__32445),
            .I(N__32278));
    InMux I__5933 (
            .O(N__32444),
            .I(N__32261));
    InMux I__5932 (
            .O(N__32443),
            .I(N__32261));
    InMux I__5931 (
            .O(N__32440),
            .I(N__32261));
    InMux I__5930 (
            .O(N__32439),
            .I(N__32261));
    InMux I__5929 (
            .O(N__32436),
            .I(N__32261));
    InMux I__5928 (
            .O(N__32435),
            .I(N__32261));
    InMux I__5927 (
            .O(N__32432),
            .I(N__32261));
    InMux I__5926 (
            .O(N__32431),
            .I(N__32261));
    Span4Mux_h I__5925 (
            .O(N__32428),
            .I(N__32250));
    Span4Mux_h I__5924 (
            .O(N__32423),
            .I(N__32250));
    LocalMux I__5923 (
            .O(N__32410),
            .I(N__32250));
    LocalMux I__5922 (
            .O(N__32395),
            .I(N__32250));
    LocalMux I__5921 (
            .O(N__32378),
            .I(N__32250));
    InMux I__5920 (
            .O(N__32375),
            .I(N__32233));
    InMux I__5919 (
            .O(N__32374),
            .I(N__32233));
    InMux I__5918 (
            .O(N__32371),
            .I(N__32233));
    InMux I__5917 (
            .O(N__32370),
            .I(N__32233));
    InMux I__5916 (
            .O(N__32367),
            .I(N__32233));
    InMux I__5915 (
            .O(N__32366),
            .I(N__32233));
    InMux I__5914 (
            .O(N__32363),
            .I(N__32233));
    InMux I__5913 (
            .O(N__32362),
            .I(N__32233));
    InMux I__5912 (
            .O(N__32359),
            .I(N__32216));
    InMux I__5911 (
            .O(N__32358),
            .I(N__32216));
    InMux I__5910 (
            .O(N__32355),
            .I(N__32216));
    InMux I__5909 (
            .O(N__32354),
            .I(N__32216));
    InMux I__5908 (
            .O(N__32351),
            .I(N__32216));
    InMux I__5907 (
            .O(N__32350),
            .I(N__32216));
    InMux I__5906 (
            .O(N__32347),
            .I(N__32216));
    InMux I__5905 (
            .O(N__32346),
            .I(N__32216));
    InMux I__5904 (
            .O(N__32343),
            .I(N__32199));
    InMux I__5903 (
            .O(N__32342),
            .I(N__32199));
    InMux I__5902 (
            .O(N__32339),
            .I(N__32199));
    InMux I__5901 (
            .O(N__32338),
            .I(N__32199));
    InMux I__5900 (
            .O(N__32335),
            .I(N__32199));
    InMux I__5899 (
            .O(N__32334),
            .I(N__32199));
    InMux I__5898 (
            .O(N__32331),
            .I(N__32199));
    InMux I__5897 (
            .O(N__32330),
            .I(N__32199));
    InMux I__5896 (
            .O(N__32327),
            .I(N__32186));
    InMux I__5895 (
            .O(N__32326),
            .I(N__32186));
    InMux I__5894 (
            .O(N__32323),
            .I(N__32186));
    InMux I__5893 (
            .O(N__32322),
            .I(N__32186));
    InMux I__5892 (
            .O(N__32319),
            .I(N__32186));
    InMux I__5891 (
            .O(N__32318),
            .I(N__32186));
    Span4Mux_v I__5890 (
            .O(N__32309),
            .I(N__32183));
    Odrv4 I__5889 (
            .O(N__32306),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__5888 (
            .O(N__32303),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5887 (
            .O(N__32288),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5886 (
            .O(N__32281),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5885 (
            .O(N__32278),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5884 (
            .O(N__32261),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__5883 (
            .O(N__32250),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5882 (
            .O(N__32233),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5881 (
            .O(N__32216),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5880 (
            .O(N__32199),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__5879 (
            .O(N__32186),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__5878 (
            .O(N__32183),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    InMux I__5877 (
            .O(N__32158),
            .I(N__32148));
    InMux I__5876 (
            .O(N__32157),
            .I(N__32148));
    InMux I__5875 (
            .O(N__32156),
            .I(N__32148));
    CascadeMux I__5874 (
            .O(N__32155),
            .I(N__32143));
    LocalMux I__5873 (
            .O(N__32148),
            .I(N__32129));
    InMux I__5872 (
            .O(N__32147),
            .I(N__32125));
    InMux I__5871 (
            .O(N__32146),
            .I(N__32096));
    InMux I__5870 (
            .O(N__32143),
            .I(N__32096));
    InMux I__5869 (
            .O(N__32142),
            .I(N__32096));
    InMux I__5868 (
            .O(N__32141),
            .I(N__32096));
    InMux I__5867 (
            .O(N__32140),
            .I(N__32096));
    CascadeMux I__5866 (
            .O(N__32139),
            .I(N__32093));
    InMux I__5865 (
            .O(N__32138),
            .I(N__32083));
    InMux I__5864 (
            .O(N__32137),
            .I(N__32070));
    InMux I__5863 (
            .O(N__32136),
            .I(N__32070));
    InMux I__5862 (
            .O(N__32135),
            .I(N__32070));
    InMux I__5861 (
            .O(N__32134),
            .I(N__32070));
    InMux I__5860 (
            .O(N__32133),
            .I(N__32070));
    InMux I__5859 (
            .O(N__32132),
            .I(N__32070));
    Span4Mux_v I__5858 (
            .O(N__32129),
            .I(N__32067));
    InMux I__5857 (
            .O(N__32128),
            .I(N__32064));
    LocalMux I__5856 (
            .O(N__32125),
            .I(N__32061));
    InMux I__5855 (
            .O(N__32124),
            .I(N__32050));
    InMux I__5854 (
            .O(N__32123),
            .I(N__32050));
    InMux I__5853 (
            .O(N__32122),
            .I(N__32050));
    InMux I__5852 (
            .O(N__32121),
            .I(N__32050));
    InMux I__5851 (
            .O(N__32120),
            .I(N__32050));
    InMux I__5850 (
            .O(N__32119),
            .I(N__32037));
    InMux I__5849 (
            .O(N__32118),
            .I(N__32037));
    InMux I__5848 (
            .O(N__32117),
            .I(N__32037));
    InMux I__5847 (
            .O(N__32116),
            .I(N__32037));
    InMux I__5846 (
            .O(N__32115),
            .I(N__32037));
    InMux I__5845 (
            .O(N__32114),
            .I(N__32037));
    InMux I__5844 (
            .O(N__32113),
            .I(N__32026));
    InMux I__5843 (
            .O(N__32112),
            .I(N__32026));
    InMux I__5842 (
            .O(N__32111),
            .I(N__32026));
    InMux I__5841 (
            .O(N__32110),
            .I(N__32026));
    InMux I__5840 (
            .O(N__32109),
            .I(N__32026));
    InMux I__5839 (
            .O(N__32108),
            .I(N__32022));
    CascadeMux I__5838 (
            .O(N__32107),
            .I(N__32019));
    LocalMux I__5837 (
            .O(N__32096),
            .I(N__32011));
    InMux I__5836 (
            .O(N__32093),
            .I(N__31994));
    InMux I__5835 (
            .O(N__32092),
            .I(N__31994));
    InMux I__5834 (
            .O(N__32091),
            .I(N__31994));
    InMux I__5833 (
            .O(N__32090),
            .I(N__31994));
    InMux I__5832 (
            .O(N__32089),
            .I(N__31994));
    InMux I__5831 (
            .O(N__32088),
            .I(N__31994));
    InMux I__5830 (
            .O(N__32087),
            .I(N__31994));
    InMux I__5829 (
            .O(N__32086),
            .I(N__31994));
    LocalMux I__5828 (
            .O(N__32083),
            .I(N__31982));
    LocalMux I__5827 (
            .O(N__32070),
            .I(N__31977));
    Span4Mux_h I__5826 (
            .O(N__32067),
            .I(N__31977));
    LocalMux I__5825 (
            .O(N__32064),
            .I(N__31968));
    Span4Mux_v I__5824 (
            .O(N__32061),
            .I(N__31968));
    LocalMux I__5823 (
            .O(N__32050),
            .I(N__31968));
    LocalMux I__5822 (
            .O(N__32037),
            .I(N__31968));
    LocalMux I__5821 (
            .O(N__32026),
            .I(N__31965));
    CascadeMux I__5820 (
            .O(N__32025),
            .I(N__31953));
    LocalMux I__5819 (
            .O(N__32022),
            .I(N__31946));
    InMux I__5818 (
            .O(N__32019),
            .I(N__31933));
    InMux I__5817 (
            .O(N__32018),
            .I(N__31933));
    InMux I__5816 (
            .O(N__32017),
            .I(N__31933));
    InMux I__5815 (
            .O(N__32016),
            .I(N__31933));
    InMux I__5814 (
            .O(N__32015),
            .I(N__31933));
    InMux I__5813 (
            .O(N__32014),
            .I(N__31933));
    Span4Mux_v I__5812 (
            .O(N__32011),
            .I(N__31928));
    LocalMux I__5811 (
            .O(N__31994),
            .I(N__31928));
    InMux I__5810 (
            .O(N__31993),
            .I(N__31913));
    InMux I__5809 (
            .O(N__31992),
            .I(N__31913));
    InMux I__5808 (
            .O(N__31991),
            .I(N__31913));
    InMux I__5807 (
            .O(N__31990),
            .I(N__31913));
    InMux I__5806 (
            .O(N__31989),
            .I(N__31913));
    InMux I__5805 (
            .O(N__31988),
            .I(N__31913));
    InMux I__5804 (
            .O(N__31987),
            .I(N__31913));
    InMux I__5803 (
            .O(N__31986),
            .I(N__31908));
    InMux I__5802 (
            .O(N__31985),
            .I(N__31908));
    Span12Mux_s11_h I__5801 (
            .O(N__31982),
            .I(N__31905));
    Span4Mux_v I__5800 (
            .O(N__31977),
            .I(N__31902));
    Span4Mux_v I__5799 (
            .O(N__31968),
            .I(N__31897));
    Span4Mux_v I__5798 (
            .O(N__31965),
            .I(N__31897));
    InMux I__5797 (
            .O(N__31964),
            .I(N__31882));
    InMux I__5796 (
            .O(N__31963),
            .I(N__31882));
    InMux I__5795 (
            .O(N__31962),
            .I(N__31882));
    InMux I__5794 (
            .O(N__31961),
            .I(N__31882));
    InMux I__5793 (
            .O(N__31960),
            .I(N__31882));
    InMux I__5792 (
            .O(N__31959),
            .I(N__31882));
    InMux I__5791 (
            .O(N__31958),
            .I(N__31882));
    InMux I__5790 (
            .O(N__31957),
            .I(N__31879));
    InMux I__5789 (
            .O(N__31956),
            .I(N__31866));
    InMux I__5788 (
            .O(N__31953),
            .I(N__31866));
    InMux I__5787 (
            .O(N__31952),
            .I(N__31866));
    InMux I__5786 (
            .O(N__31951),
            .I(N__31866));
    InMux I__5785 (
            .O(N__31950),
            .I(N__31866));
    InMux I__5784 (
            .O(N__31949),
            .I(N__31866));
    Span4Mux_h I__5783 (
            .O(N__31946),
            .I(N__31859));
    LocalMux I__5782 (
            .O(N__31933),
            .I(N__31859));
    Span4Mux_h I__5781 (
            .O(N__31928),
            .I(N__31859));
    LocalMux I__5780 (
            .O(N__31913),
            .I(N__31854));
    LocalMux I__5779 (
            .O(N__31908),
            .I(N__31854));
    Odrv12 I__5778 (
            .O(N__31905),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5777 (
            .O(N__31902),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5776 (
            .O(N__31897),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__5775 (
            .O(N__31882),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__5774 (
            .O(N__31879),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__5773 (
            .O(N__31866),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__5772 (
            .O(N__31859),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__5771 (
            .O(N__31854),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__5770 (
            .O(N__31837),
            .I(N__31834));
    InMux I__5769 (
            .O(N__31834),
            .I(N__31831));
    LocalMux I__5768 (
            .O(N__31831),
            .I(N__31826));
    InMux I__5767 (
            .O(N__31830),
            .I(N__31823));
    InMux I__5766 (
            .O(N__31829),
            .I(N__31820));
    Span12Mux_h I__5765 (
            .O(N__31826),
            .I(N__31817));
    LocalMux I__5764 (
            .O(N__31823),
            .I(N__31814));
    LocalMux I__5763 (
            .O(N__31820),
            .I(N__31811));
    Odrv12 I__5762 (
            .O(N__31817),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv12 I__5761 (
            .O(N__31814),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__5760 (
            .O(N__31811),
            .I(\current_shift_inst.un4_control_input1_20 ));
    CascadeMux I__5759 (
            .O(N__31804),
            .I(N__31800));
    InMux I__5758 (
            .O(N__31803),
            .I(N__31797));
    InMux I__5757 (
            .O(N__31800),
            .I(N__31794));
    LocalMux I__5756 (
            .O(N__31797),
            .I(N__31789));
    LocalMux I__5755 (
            .O(N__31794),
            .I(N__31789));
    Span4Mux_v I__5754 (
            .O(N__31789),
            .I(N__31785));
    CascadeMux I__5753 (
            .O(N__31788),
            .I(N__31782));
    Span4Mux_h I__5752 (
            .O(N__31785),
            .I(N__31778));
    InMux I__5751 (
            .O(N__31782),
            .I(N__31775));
    InMux I__5750 (
            .O(N__31781),
            .I(N__31772));
    Span4Mux_h I__5749 (
            .O(N__31778),
            .I(N__31767));
    LocalMux I__5748 (
            .O(N__31775),
            .I(N__31767));
    LocalMux I__5747 (
            .O(N__31772),
            .I(N__31764));
    Odrv4 I__5746 (
            .O(N__31767),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__5745 (
            .O(N__31764),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__5744 (
            .O(N__31759),
            .I(N__31756));
    LocalMux I__5743 (
            .O(N__31756),
            .I(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ));
    CascadeMux I__5742 (
            .O(N__31753),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_ ));
    CascadeMux I__5741 (
            .O(N__31750),
            .I(elapsed_time_ns_1_RNIRB3CP1_0_3_cascade_));
    InMux I__5740 (
            .O(N__31747),
            .I(N__31744));
    LocalMux I__5739 (
            .O(N__31744),
            .I(N__31741));
    Span4Mux_v I__5738 (
            .O(N__31741),
            .I(N__31738));
    Odrv4 I__5737 (
            .O(N__31738),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__5736 (
            .O(N__31735),
            .I(N__31732));
    LocalMux I__5735 (
            .O(N__31732),
            .I(N__31729));
    Odrv4 I__5734 (
            .O(N__31729),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__5733 (
            .O(N__31726),
            .I(N__31723));
    InMux I__5732 (
            .O(N__31723),
            .I(N__31720));
    LocalMux I__5731 (
            .O(N__31720),
            .I(N__31717));
    Odrv4 I__5730 (
            .O(N__31717),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__5729 (
            .O(N__31714),
            .I(N__31711));
    InMux I__5728 (
            .O(N__31711),
            .I(N__31708));
    LocalMux I__5727 (
            .O(N__31708),
            .I(N__31705));
    Odrv4 I__5726 (
            .O(N__31705),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__5725 (
            .O(N__31702),
            .I(N__31699));
    LocalMux I__5724 (
            .O(N__31699),
            .I(N__31696));
    Odrv4 I__5723 (
            .O(N__31696),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__5722 (
            .O(N__31693),
            .I(N__31690));
    LocalMux I__5721 (
            .O(N__31690),
            .I(N__31687));
    Span4Mux_v I__5720 (
            .O(N__31687),
            .I(N__31684));
    Odrv4 I__5719 (
            .O(N__31684),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__5718 (
            .O(N__31681),
            .I(N__31678));
    LocalMux I__5717 (
            .O(N__31678),
            .I(N__31675));
    Odrv4 I__5716 (
            .O(N__31675),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__5715 (
            .O(N__31672),
            .I(N__31669));
    LocalMux I__5714 (
            .O(N__31669),
            .I(N__31666));
    Span4Mux_h I__5713 (
            .O(N__31666),
            .I(N__31663));
    Span4Mux_v I__5712 (
            .O(N__31663),
            .I(N__31660));
    Odrv4 I__5711 (
            .O(N__31660),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__5710 (
            .O(N__31657),
            .I(N__31654));
    LocalMux I__5709 (
            .O(N__31654),
            .I(N__31649));
    InMux I__5708 (
            .O(N__31653),
            .I(N__31646));
    InMux I__5707 (
            .O(N__31652),
            .I(N__31643));
    Span4Mux_h I__5706 (
            .O(N__31649),
            .I(N__31639));
    LocalMux I__5705 (
            .O(N__31646),
            .I(N__31636));
    LocalMux I__5704 (
            .O(N__31643),
            .I(N__31633));
    InMux I__5703 (
            .O(N__31642),
            .I(N__31630));
    Span4Mux_v I__5702 (
            .O(N__31639),
            .I(N__31627));
    Span4Mux_h I__5701 (
            .O(N__31636),
            .I(N__31624));
    Span12Mux_h I__5700 (
            .O(N__31633),
            .I(N__31619));
    LocalMux I__5699 (
            .O(N__31630),
            .I(N__31619));
    Odrv4 I__5698 (
            .O(N__31627),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__5697 (
            .O(N__31624),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv12 I__5696 (
            .O(N__31619),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    CascadeMux I__5695 (
            .O(N__31612),
            .I(N__31609));
    InMux I__5694 (
            .O(N__31609),
            .I(N__31605));
    CascadeMux I__5693 (
            .O(N__31608),
            .I(N__31602));
    LocalMux I__5692 (
            .O(N__31605),
            .I(N__31599));
    InMux I__5691 (
            .O(N__31602),
            .I(N__31596));
    Span4Mux_v I__5690 (
            .O(N__31599),
            .I(N__31590));
    LocalMux I__5689 (
            .O(N__31596),
            .I(N__31590));
    InMux I__5688 (
            .O(N__31595),
            .I(N__31587));
    Span4Mux_h I__5687 (
            .O(N__31590),
            .I(N__31584));
    LocalMux I__5686 (
            .O(N__31587),
            .I(N__31581));
    Odrv4 I__5685 (
            .O(N__31584),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv12 I__5684 (
            .O(N__31581),
            .I(\current_shift_inst.un4_control_input1_25 ));
    CascadeMux I__5683 (
            .O(N__31576),
            .I(N__31573));
    InMux I__5682 (
            .O(N__31573),
            .I(N__31570));
    LocalMux I__5681 (
            .O(N__31570),
            .I(N__31567));
    Odrv4 I__5680 (
            .O(N__31567),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    CascadeMux I__5679 (
            .O(N__31564),
            .I(N__31560));
    CascadeMux I__5678 (
            .O(N__31563),
            .I(N__31557));
    InMux I__5677 (
            .O(N__31560),
            .I(N__31554));
    InMux I__5676 (
            .O(N__31557),
            .I(N__31551));
    LocalMux I__5675 (
            .O(N__31554),
            .I(N__31548));
    LocalMux I__5674 (
            .O(N__31551),
            .I(N__31545));
    Span4Mux_h I__5673 (
            .O(N__31548),
            .I(N__31540));
    Span4Mux_h I__5672 (
            .O(N__31545),
            .I(N__31537));
    InMux I__5671 (
            .O(N__31544),
            .I(N__31534));
    InMux I__5670 (
            .O(N__31543),
            .I(N__31531));
    Span4Mux_v I__5669 (
            .O(N__31540),
            .I(N__31528));
    Span4Mux_h I__5668 (
            .O(N__31537),
            .I(N__31521));
    LocalMux I__5667 (
            .O(N__31534),
            .I(N__31521));
    LocalMux I__5666 (
            .O(N__31531),
            .I(N__31521));
    Odrv4 I__5665 (
            .O(N__31528),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__5664 (
            .O(N__31521),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__5663 (
            .O(N__31516),
            .I(N__31513));
    LocalMux I__5662 (
            .O(N__31513),
            .I(N__31509));
    InMux I__5661 (
            .O(N__31512),
            .I(N__31505));
    Span4Mux_h I__5660 (
            .O(N__31509),
            .I(N__31502));
    InMux I__5659 (
            .O(N__31508),
            .I(N__31499));
    LocalMux I__5658 (
            .O(N__31505),
            .I(N__31496));
    Odrv4 I__5657 (
            .O(N__31502),
            .I(\current_shift_inst.un4_control_input1_24 ));
    LocalMux I__5656 (
            .O(N__31499),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv12 I__5655 (
            .O(N__31496),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__5654 (
            .O(N__31489),
            .I(N__31486));
    LocalMux I__5653 (
            .O(N__31486),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__5652 (
            .O(N__31483),
            .I(N__31480));
    LocalMux I__5651 (
            .O(N__31480),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__5650 (
            .O(N__31477),
            .I(N__31474));
    LocalMux I__5649 (
            .O(N__31474),
            .I(N__31471));
    Span4Mux_v I__5648 (
            .O(N__31471),
            .I(N__31468));
    Odrv4 I__5647 (
            .O(N__31468),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__5646 (
            .O(N__31465),
            .I(N__31462));
    LocalMux I__5645 (
            .O(N__31462),
            .I(N__31459));
    Odrv12 I__5644 (
            .O(N__31459),
            .I(\current_shift_inst.control_input_axb_9 ));
    CascadeMux I__5643 (
            .O(N__31456),
            .I(N__31453));
    InMux I__5642 (
            .O(N__31453),
            .I(N__31450));
    LocalMux I__5641 (
            .O(N__31450),
            .I(N__31446));
    InMux I__5640 (
            .O(N__31449),
            .I(N__31443));
    Span4Mux_v I__5639 (
            .O(N__31446),
            .I(N__31439));
    LocalMux I__5638 (
            .O(N__31443),
            .I(N__31436));
    InMux I__5637 (
            .O(N__31442),
            .I(N__31433));
    Span4Mux_h I__5636 (
            .O(N__31439),
            .I(N__31428));
    Span4Mux_v I__5635 (
            .O(N__31436),
            .I(N__31428));
    LocalMux I__5634 (
            .O(N__31433),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__5633 (
            .O(N__31428),
            .I(\current_shift_inst.un4_control_input1_11 ));
    CascadeMux I__5632 (
            .O(N__31423),
            .I(N__31420));
    InMux I__5631 (
            .O(N__31420),
            .I(N__31416));
    InMux I__5630 (
            .O(N__31419),
            .I(N__31413));
    LocalMux I__5629 (
            .O(N__31416),
            .I(N__31410));
    LocalMux I__5628 (
            .O(N__31413),
            .I(N__31407));
    Span4Mux_h I__5627 (
            .O(N__31410),
            .I(N__31403));
    Span4Mux_v I__5626 (
            .O(N__31407),
            .I(N__31400));
    InMux I__5625 (
            .O(N__31406),
            .I(N__31397));
    Span4Mux_v I__5624 (
            .O(N__31403),
            .I(N__31393));
    Span4Mux_h I__5623 (
            .O(N__31400),
            .I(N__31388));
    LocalMux I__5622 (
            .O(N__31397),
            .I(N__31388));
    InMux I__5621 (
            .O(N__31396),
            .I(N__31385));
    Odrv4 I__5620 (
            .O(N__31393),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__5619 (
            .O(N__31388),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__5618 (
            .O(N__31385),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    CascadeMux I__5617 (
            .O(N__31378),
            .I(N__31375));
    InMux I__5616 (
            .O(N__31375),
            .I(N__31372));
    LocalMux I__5615 (
            .O(N__31372),
            .I(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ));
    CascadeMux I__5614 (
            .O(N__31369),
            .I(N__31365));
    CascadeMux I__5613 (
            .O(N__31368),
            .I(N__31362));
    InMux I__5612 (
            .O(N__31365),
            .I(N__31359));
    InMux I__5611 (
            .O(N__31362),
            .I(N__31356));
    LocalMux I__5610 (
            .O(N__31359),
            .I(N__31353));
    LocalMux I__5609 (
            .O(N__31356),
            .I(N__31348));
    Span4Mux_h I__5608 (
            .O(N__31353),
            .I(N__31345));
    InMux I__5607 (
            .O(N__31352),
            .I(N__31342));
    InMux I__5606 (
            .O(N__31351),
            .I(N__31339));
    Span4Mux_v I__5605 (
            .O(N__31348),
            .I(N__31336));
    Span4Mux_v I__5604 (
            .O(N__31345),
            .I(N__31331));
    LocalMux I__5603 (
            .O(N__31342),
            .I(N__31331));
    LocalMux I__5602 (
            .O(N__31339),
            .I(N__31328));
    Span4Mux_h I__5601 (
            .O(N__31336),
            .I(N__31325));
    Span4Mux_h I__5600 (
            .O(N__31331),
            .I(N__31322));
    Span4Mux_v I__5599 (
            .O(N__31328),
            .I(N__31319));
    Odrv4 I__5598 (
            .O(N__31325),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__5597 (
            .O(N__31322),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__5596 (
            .O(N__31319),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__5595 (
            .O(N__31312),
            .I(N__31308));
    InMux I__5594 (
            .O(N__31311),
            .I(N__31305));
    LocalMux I__5593 (
            .O(N__31308),
            .I(N__31302));
    LocalMux I__5592 (
            .O(N__31305),
            .I(N__31298));
    Span4Mux_h I__5591 (
            .O(N__31302),
            .I(N__31295));
    InMux I__5590 (
            .O(N__31301),
            .I(N__31292));
    Span4Mux_v I__5589 (
            .O(N__31298),
            .I(N__31289));
    Odrv4 I__5588 (
            .O(N__31295),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__5587 (
            .O(N__31292),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__5586 (
            .O(N__31289),
            .I(\current_shift_inst.un4_control_input1_15 ));
    CascadeMux I__5585 (
            .O(N__31282),
            .I(N__31279));
    InMux I__5584 (
            .O(N__31279),
            .I(N__31276));
    LocalMux I__5583 (
            .O(N__31276),
            .I(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ));
    CascadeMux I__5582 (
            .O(N__31273),
            .I(N__31270));
    InMux I__5581 (
            .O(N__31270),
            .I(N__31267));
    LocalMux I__5580 (
            .O(N__31267),
            .I(N__31263));
    InMux I__5579 (
            .O(N__31266),
            .I(N__31259));
    Span4Mux_h I__5578 (
            .O(N__31263),
            .I(N__31256));
    InMux I__5577 (
            .O(N__31262),
            .I(N__31253));
    LocalMux I__5576 (
            .O(N__31259),
            .I(N__31250));
    Odrv4 I__5575 (
            .O(N__31256),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__5574 (
            .O(N__31253),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__5573 (
            .O(N__31250),
            .I(\current_shift_inst.un4_control_input1_23 ));
    CascadeMux I__5572 (
            .O(N__31243),
            .I(N__31240));
    InMux I__5571 (
            .O(N__31240),
            .I(N__31236));
    InMux I__5570 (
            .O(N__31239),
            .I(N__31233));
    LocalMux I__5569 (
            .O(N__31236),
            .I(N__31229));
    LocalMux I__5568 (
            .O(N__31233),
            .I(N__31225));
    InMux I__5567 (
            .O(N__31232),
            .I(N__31222));
    Span4Mux_h I__5566 (
            .O(N__31229),
            .I(N__31219));
    InMux I__5565 (
            .O(N__31228),
            .I(N__31216));
    Span4Mux_h I__5564 (
            .O(N__31225),
            .I(N__31211));
    LocalMux I__5563 (
            .O(N__31222),
            .I(N__31211));
    Span4Mux_v I__5562 (
            .O(N__31219),
            .I(N__31208));
    LocalMux I__5561 (
            .O(N__31216),
            .I(N__31203));
    Span4Mux_h I__5560 (
            .O(N__31211),
            .I(N__31203));
    Odrv4 I__5559 (
            .O(N__31208),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__5558 (
            .O(N__31203),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    CascadeMux I__5557 (
            .O(N__31198),
            .I(N__31195));
    InMux I__5556 (
            .O(N__31195),
            .I(N__31192));
    LocalMux I__5555 (
            .O(N__31192),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    CascadeMux I__5554 (
            .O(N__31189),
            .I(N__31186));
    InMux I__5553 (
            .O(N__31186),
            .I(N__31183));
    LocalMux I__5552 (
            .O(N__31183),
            .I(N__31179));
    InMux I__5551 (
            .O(N__31182),
            .I(N__31176));
    Span4Mux_v I__5550 (
            .O(N__31179),
            .I(N__31173));
    LocalMux I__5549 (
            .O(N__31176),
            .I(N__31170));
    Span4Mux_v I__5548 (
            .O(N__31173),
            .I(N__31165));
    Span4Mux_h I__5547 (
            .O(N__31170),
            .I(N__31162));
    InMux I__5546 (
            .O(N__31169),
            .I(N__31159));
    InMux I__5545 (
            .O(N__31168),
            .I(N__31156));
    Span4Mux_h I__5544 (
            .O(N__31165),
            .I(N__31153));
    Span4Mux_h I__5543 (
            .O(N__31162),
            .I(N__31150));
    LocalMux I__5542 (
            .O(N__31159),
            .I(N__31145));
    LocalMux I__5541 (
            .O(N__31156),
            .I(N__31145));
    Odrv4 I__5540 (
            .O(N__31153),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__5539 (
            .O(N__31150),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv12 I__5538 (
            .O(N__31145),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__5537 (
            .O(N__31138),
            .I(N__31134));
    InMux I__5536 (
            .O(N__31137),
            .I(N__31131));
    LocalMux I__5535 (
            .O(N__31134),
            .I(N__31127));
    LocalMux I__5534 (
            .O(N__31131),
            .I(N__31124));
    InMux I__5533 (
            .O(N__31130),
            .I(N__31121));
    Span4Mux_h I__5532 (
            .O(N__31127),
            .I(N__31116));
    Span4Mux_v I__5531 (
            .O(N__31124),
            .I(N__31116));
    LocalMux I__5530 (
            .O(N__31121),
            .I(\current_shift_inst.un4_control_input1_21 ));
    Odrv4 I__5529 (
            .O(N__31116),
            .I(\current_shift_inst.un4_control_input1_21 ));
    CascadeMux I__5528 (
            .O(N__31111),
            .I(N__31108));
    InMux I__5527 (
            .O(N__31108),
            .I(N__31105));
    LocalMux I__5526 (
            .O(N__31105),
            .I(N__31102));
    Odrv12 I__5525 (
            .O(N__31102),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    CascadeMux I__5524 (
            .O(N__31099),
            .I(N__31096));
    InMux I__5523 (
            .O(N__31096),
            .I(N__31092));
    CascadeMux I__5522 (
            .O(N__31095),
            .I(N__31089));
    LocalMux I__5521 (
            .O(N__31092),
            .I(N__31085));
    InMux I__5520 (
            .O(N__31089),
            .I(N__31082));
    InMux I__5519 (
            .O(N__31088),
            .I(N__31079));
    Span4Mux_h I__5518 (
            .O(N__31085),
            .I(N__31076));
    LocalMux I__5517 (
            .O(N__31082),
            .I(N__31073));
    LocalMux I__5516 (
            .O(N__31079),
            .I(N__31070));
    Odrv4 I__5515 (
            .O(N__31076),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv12 I__5514 (
            .O(N__31073),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv12 I__5513 (
            .O(N__31070),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__5512 (
            .O(N__31063),
            .I(N__31060));
    LocalMux I__5511 (
            .O(N__31060),
            .I(N__31055));
    InMux I__5510 (
            .O(N__31059),
            .I(N__31052));
    InMux I__5509 (
            .O(N__31058),
            .I(N__31049));
    Span4Mux_v I__5508 (
            .O(N__31055),
            .I(N__31043));
    LocalMux I__5507 (
            .O(N__31052),
            .I(N__31043));
    LocalMux I__5506 (
            .O(N__31049),
            .I(N__31040));
    InMux I__5505 (
            .O(N__31048),
            .I(N__31037));
    Span4Mux_h I__5504 (
            .O(N__31043),
            .I(N__31034));
    Span12Mux_h I__5503 (
            .O(N__31040),
            .I(N__31029));
    LocalMux I__5502 (
            .O(N__31037),
            .I(N__31029));
    Odrv4 I__5501 (
            .O(N__31034),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv12 I__5500 (
            .O(N__31029),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__5499 (
            .O(N__31024),
            .I(N__31021));
    LocalMux I__5498 (
            .O(N__31021),
            .I(N__31018));
    Odrv12 I__5497 (
            .O(N__31018),
            .I(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ));
    CascadeMux I__5496 (
            .O(N__31015),
            .I(N__31011));
    CascadeMux I__5495 (
            .O(N__31014),
            .I(N__31008));
    InMux I__5494 (
            .O(N__31011),
            .I(N__31005));
    InMux I__5493 (
            .O(N__31008),
            .I(N__31002));
    LocalMux I__5492 (
            .O(N__31005),
            .I(N__30998));
    LocalMux I__5491 (
            .O(N__31002),
            .I(N__30995));
    InMux I__5490 (
            .O(N__31001),
            .I(N__30992));
    Span4Mux_h I__5489 (
            .O(N__30998),
            .I(N__30985));
    Span4Mux_v I__5488 (
            .O(N__30995),
            .I(N__30985));
    LocalMux I__5487 (
            .O(N__30992),
            .I(N__30985));
    Span4Mux_h I__5486 (
            .O(N__30985),
            .I(N__30982));
    Span4Mux_v I__5485 (
            .O(N__30982),
            .I(N__30978));
    InMux I__5484 (
            .O(N__30981),
            .I(N__30975));
    Odrv4 I__5483 (
            .O(N__30978),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__5482 (
            .O(N__30975),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__5481 (
            .O(N__30970),
            .I(N__30967));
    LocalMux I__5480 (
            .O(N__30967),
            .I(N__30964));
    Span4Mux_h I__5479 (
            .O(N__30964),
            .I(N__30959));
    InMux I__5478 (
            .O(N__30963),
            .I(N__30956));
    InMux I__5477 (
            .O(N__30962),
            .I(N__30953));
    Odrv4 I__5476 (
            .O(N__30959),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__5475 (
            .O(N__30956),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__5474 (
            .O(N__30953),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__5473 (
            .O(N__30946),
            .I(N__30943));
    LocalMux I__5472 (
            .O(N__30943),
            .I(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ));
    CascadeMux I__5471 (
            .O(N__30940),
            .I(N__30936));
    CascadeMux I__5470 (
            .O(N__30939),
            .I(N__30933));
    InMux I__5469 (
            .O(N__30936),
            .I(N__30930));
    InMux I__5468 (
            .O(N__30933),
            .I(N__30927));
    LocalMux I__5467 (
            .O(N__30930),
            .I(N__30924));
    LocalMux I__5466 (
            .O(N__30927),
            .I(N__30920));
    Span4Mux_v I__5465 (
            .O(N__30924),
            .I(N__30916));
    InMux I__5464 (
            .O(N__30923),
            .I(N__30913));
    Span4Mux_h I__5463 (
            .O(N__30920),
            .I(N__30910));
    InMux I__5462 (
            .O(N__30919),
            .I(N__30907));
    Span4Mux_h I__5461 (
            .O(N__30916),
            .I(N__30902));
    LocalMux I__5460 (
            .O(N__30913),
            .I(N__30902));
    Sp12to4 I__5459 (
            .O(N__30910),
            .I(N__30897));
    LocalMux I__5458 (
            .O(N__30907),
            .I(N__30897));
    Odrv4 I__5457 (
            .O(N__30902),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv12 I__5456 (
            .O(N__30897),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__5455 (
            .O(N__30892),
            .I(N__30889));
    LocalMux I__5454 (
            .O(N__30889),
            .I(N__30885));
    InMux I__5453 (
            .O(N__30888),
            .I(N__30881));
    Span4Mux_v I__5452 (
            .O(N__30885),
            .I(N__30878));
    InMux I__5451 (
            .O(N__30884),
            .I(N__30875));
    LocalMux I__5450 (
            .O(N__30881),
            .I(N__30872));
    Odrv4 I__5449 (
            .O(N__30878),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__5448 (
            .O(N__30875),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv12 I__5447 (
            .O(N__30872),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__5446 (
            .O(N__30865),
            .I(N__30862));
    LocalMux I__5445 (
            .O(N__30862),
            .I(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ));
    InMux I__5444 (
            .O(N__30859),
            .I(N__30856));
    LocalMux I__5443 (
            .O(N__30856),
            .I(N__30853));
    Odrv4 I__5442 (
            .O(N__30853),
            .I(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ));
    CascadeMux I__5441 (
            .O(N__30850),
            .I(N__30846));
    CascadeMux I__5440 (
            .O(N__30849),
            .I(N__30843));
    InMux I__5439 (
            .O(N__30846),
            .I(N__30840));
    InMux I__5438 (
            .O(N__30843),
            .I(N__30837));
    LocalMux I__5437 (
            .O(N__30840),
            .I(N__30834));
    LocalMux I__5436 (
            .O(N__30837),
            .I(N__30831));
    Span4Mux_h I__5435 (
            .O(N__30834),
            .I(N__30826));
    Span4Mux_v I__5434 (
            .O(N__30831),
            .I(N__30823));
    InMux I__5433 (
            .O(N__30830),
            .I(N__30820));
    InMux I__5432 (
            .O(N__30829),
            .I(N__30817));
    Span4Mux_v I__5431 (
            .O(N__30826),
            .I(N__30814));
    Span4Mux_h I__5430 (
            .O(N__30823),
            .I(N__30809));
    LocalMux I__5429 (
            .O(N__30820),
            .I(N__30809));
    LocalMux I__5428 (
            .O(N__30817),
            .I(N__30806));
    Odrv4 I__5427 (
            .O(N__30814),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__5426 (
            .O(N__30809),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv12 I__5425 (
            .O(N__30806),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__5424 (
            .O(N__30799),
            .I(N__30795));
    InMux I__5423 (
            .O(N__30798),
            .I(N__30792));
    LocalMux I__5422 (
            .O(N__30795),
            .I(N__30788));
    LocalMux I__5421 (
            .O(N__30792),
            .I(N__30785));
    InMux I__5420 (
            .O(N__30791),
            .I(N__30782));
    Span4Mux_v I__5419 (
            .O(N__30788),
            .I(N__30777));
    Span4Mux_v I__5418 (
            .O(N__30785),
            .I(N__30777));
    LocalMux I__5417 (
            .O(N__30782),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__5416 (
            .O(N__30777),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__5415 (
            .O(N__30772),
            .I(N__30769));
    LocalMux I__5414 (
            .O(N__30769),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    CascadeMux I__5413 (
            .O(N__30766),
            .I(N__30762));
    CascadeMux I__5412 (
            .O(N__30765),
            .I(N__30759));
    InMux I__5411 (
            .O(N__30762),
            .I(N__30756));
    InMux I__5410 (
            .O(N__30759),
            .I(N__30753));
    LocalMux I__5409 (
            .O(N__30756),
            .I(N__30750));
    LocalMux I__5408 (
            .O(N__30753),
            .I(N__30746));
    Span4Mux_h I__5407 (
            .O(N__30750),
            .I(N__30742));
    InMux I__5406 (
            .O(N__30749),
            .I(N__30739));
    Span4Mux_h I__5405 (
            .O(N__30746),
            .I(N__30736));
    InMux I__5404 (
            .O(N__30745),
            .I(N__30733));
    Span4Mux_h I__5403 (
            .O(N__30742),
            .I(N__30728));
    LocalMux I__5402 (
            .O(N__30739),
            .I(N__30728));
    Sp12to4 I__5401 (
            .O(N__30736),
            .I(N__30723));
    LocalMux I__5400 (
            .O(N__30733),
            .I(N__30723));
    Odrv4 I__5399 (
            .O(N__30728),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv12 I__5398 (
            .O(N__30723),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__5397 (
            .O(N__30718),
            .I(N__30715));
    LocalMux I__5396 (
            .O(N__30715),
            .I(N__30710));
    InMux I__5395 (
            .O(N__30714),
            .I(N__30707));
    InMux I__5394 (
            .O(N__30713),
            .I(N__30704));
    Span12Mux_v I__5393 (
            .O(N__30710),
            .I(N__30701));
    LocalMux I__5392 (
            .O(N__30707),
            .I(N__30698));
    LocalMux I__5391 (
            .O(N__30704),
            .I(\current_shift_inst.un4_control_input1_6 ));
    Odrv12 I__5390 (
            .O(N__30701),
            .I(\current_shift_inst.un4_control_input1_6 ));
    Odrv4 I__5389 (
            .O(N__30698),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__5388 (
            .O(N__30691),
            .I(N__30688));
    LocalMux I__5387 (
            .O(N__30688),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    CascadeMux I__5386 (
            .O(N__30685),
            .I(N__30682));
    InMux I__5385 (
            .O(N__30682),
            .I(N__30676));
    InMux I__5384 (
            .O(N__30681),
            .I(N__30676));
    LocalMux I__5383 (
            .O(N__30676),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    CascadeMux I__5382 (
            .O(N__30673),
            .I(N__30670));
    InMux I__5381 (
            .O(N__30670),
            .I(N__30661));
    InMux I__5380 (
            .O(N__30669),
            .I(N__30661));
    InMux I__5379 (
            .O(N__30668),
            .I(N__30661));
    LocalMux I__5378 (
            .O(N__30661),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__5377 (
            .O(N__30658),
            .I(N__30649));
    InMux I__5376 (
            .O(N__30657),
            .I(N__30639));
    InMux I__5375 (
            .O(N__30656),
            .I(N__30636));
    InMux I__5374 (
            .O(N__30655),
            .I(N__30631));
    InMux I__5373 (
            .O(N__30654),
            .I(N__30631));
    InMux I__5372 (
            .O(N__30653),
            .I(N__30625));
    InMux I__5371 (
            .O(N__30652),
            .I(N__30625));
    LocalMux I__5370 (
            .O(N__30649),
            .I(N__30612));
    InMux I__5369 (
            .O(N__30648),
            .I(N__30597));
    InMux I__5368 (
            .O(N__30647),
            .I(N__30597));
    InMux I__5367 (
            .O(N__30646),
            .I(N__30597));
    InMux I__5366 (
            .O(N__30645),
            .I(N__30597));
    InMux I__5365 (
            .O(N__30644),
            .I(N__30597));
    InMux I__5364 (
            .O(N__30643),
            .I(N__30597));
    InMux I__5363 (
            .O(N__30642),
            .I(N__30597));
    LocalMux I__5362 (
            .O(N__30639),
            .I(N__30592));
    LocalMux I__5361 (
            .O(N__30636),
            .I(N__30592));
    LocalMux I__5360 (
            .O(N__30631),
            .I(N__30589));
    InMux I__5359 (
            .O(N__30630),
            .I(N__30586));
    LocalMux I__5358 (
            .O(N__30625),
            .I(N__30583));
    InMux I__5357 (
            .O(N__30624),
            .I(N__30578));
    InMux I__5356 (
            .O(N__30623),
            .I(N__30578));
    InMux I__5355 (
            .O(N__30622),
            .I(N__30573));
    InMux I__5354 (
            .O(N__30621),
            .I(N__30573));
    InMux I__5353 (
            .O(N__30620),
            .I(N__30570));
    InMux I__5352 (
            .O(N__30619),
            .I(N__30559));
    InMux I__5351 (
            .O(N__30618),
            .I(N__30559));
    InMux I__5350 (
            .O(N__30617),
            .I(N__30559));
    InMux I__5349 (
            .O(N__30616),
            .I(N__30559));
    InMux I__5348 (
            .O(N__30615),
            .I(N__30559));
    Span4Mux_h I__5347 (
            .O(N__30612),
            .I(N__30552));
    LocalMux I__5346 (
            .O(N__30597),
            .I(N__30552));
    Span4Mux_v I__5345 (
            .O(N__30592),
            .I(N__30552));
    Odrv4 I__5344 (
            .O(N__30589),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__5343 (
            .O(N__30586),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__5342 (
            .O(N__30583),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__5341 (
            .O(N__30578),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__5340 (
            .O(N__30573),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__5339 (
            .O(N__30570),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__5338 (
            .O(N__30559),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__5337 (
            .O(N__30552),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    CascadeMux I__5336 (
            .O(N__30535),
            .I(N__30532));
    InMux I__5335 (
            .O(N__30532),
            .I(N__30528));
    InMux I__5334 (
            .O(N__30531),
            .I(N__30525));
    LocalMux I__5333 (
            .O(N__30528),
            .I(N__30522));
    LocalMux I__5332 (
            .O(N__30525),
            .I(N__30519));
    Span4Mux_h I__5331 (
            .O(N__30522),
            .I(N__30514));
    Span4Mux_h I__5330 (
            .O(N__30519),
            .I(N__30514));
    Span4Mux_v I__5329 (
            .O(N__30514),
            .I(N__30509));
    InMux I__5328 (
            .O(N__30513),
            .I(N__30506));
    InMux I__5327 (
            .O(N__30512),
            .I(N__30503));
    Span4Mux_h I__5326 (
            .O(N__30509),
            .I(N__30500));
    LocalMux I__5325 (
            .O(N__30506),
            .I(N__30495));
    LocalMux I__5324 (
            .O(N__30503),
            .I(N__30495));
    Odrv4 I__5323 (
            .O(N__30500),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv12 I__5322 (
            .O(N__30495),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__5321 (
            .O(N__30490),
            .I(N__30487));
    LocalMux I__5320 (
            .O(N__30487),
            .I(N__30482));
    InMux I__5319 (
            .O(N__30486),
            .I(N__30479));
    InMux I__5318 (
            .O(N__30485),
            .I(N__30476));
    Span4Mux_v I__5317 (
            .O(N__30482),
            .I(N__30473));
    LocalMux I__5316 (
            .O(N__30479),
            .I(N__30470));
    LocalMux I__5315 (
            .O(N__30476),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__5314 (
            .O(N__30473),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv12 I__5313 (
            .O(N__30470),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__5312 (
            .O(N__30463),
            .I(N__30460));
    LocalMux I__5311 (
            .O(N__30460),
            .I(N__30457));
    Span4Mux_v I__5310 (
            .O(N__30457),
            .I(N__30454));
    Odrv4 I__5309 (
            .O(N__30454),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__5308 (
            .O(N__30451),
            .I(N__30448));
    LocalMux I__5307 (
            .O(N__30448),
            .I(N__30445));
    Odrv4 I__5306 (
            .O(N__30445),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__5305 (
            .O(N__30442),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__5304 (
            .O(N__30439),
            .I(N__30436));
    LocalMux I__5303 (
            .O(N__30436),
            .I(N__30433));
    Odrv4 I__5302 (
            .O(N__30433),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__5301 (
            .O(N__30430),
            .I(bfn_12_12_0_));
    InMux I__5300 (
            .O(N__30427),
            .I(N__30424));
    LocalMux I__5299 (
            .O(N__30424),
            .I(N__30421));
    Odrv4 I__5298 (
            .O(N__30421),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__5297 (
            .O(N__30418),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__5296 (
            .O(N__30415),
            .I(N__30412));
    LocalMux I__5295 (
            .O(N__30412),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__5294 (
            .O(N__30409),
            .I(N__30406));
    LocalMux I__5293 (
            .O(N__30406),
            .I(N__30403));
    Odrv4 I__5292 (
            .O(N__30403),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__5291 (
            .O(N__30400),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__5290 (
            .O(N__30397),
            .I(N__30394));
    LocalMux I__5289 (
            .O(N__30394),
            .I(N__30391));
    Span4Mux_v I__5288 (
            .O(N__30391),
            .I(N__30388));
    Odrv4 I__5287 (
            .O(N__30388),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__5286 (
            .O(N__30385),
            .I(N__30382));
    LocalMux I__5285 (
            .O(N__30382),
            .I(N__30379));
    Odrv4 I__5284 (
            .O(N__30379),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__5283 (
            .O(N__30376),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__5282 (
            .O(N__30373),
            .I(N__30370));
    LocalMux I__5281 (
            .O(N__30370),
            .I(N__30367));
    Odrv4 I__5280 (
            .O(N__30367),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__5279 (
            .O(N__30364),
            .I(N__30361));
    LocalMux I__5278 (
            .O(N__30361),
            .I(N__30358));
    Odrv4 I__5277 (
            .O(N__30358),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__5276 (
            .O(N__30355),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__5275 (
            .O(N__30352),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__5274 (
            .O(N__30349),
            .I(N__30346));
    LocalMux I__5273 (
            .O(N__30346),
            .I(N__30343));
    Odrv4 I__5272 (
            .O(N__30343),
            .I(\current_shift_inst.control_input_31 ));
    CascadeMux I__5271 (
            .O(N__30340),
            .I(\current_shift_inst.control_input_31_cascade_ ));
    InMux I__5270 (
            .O(N__30337),
            .I(N__30334));
    LocalMux I__5269 (
            .O(N__30334),
            .I(N__30331));
    Odrv4 I__5268 (
            .O(N__30331),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__5267 (
            .O(N__30328),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    CascadeMux I__5266 (
            .O(N__30325),
            .I(N__30322));
    InMux I__5265 (
            .O(N__30322),
            .I(N__30319));
    LocalMux I__5264 (
            .O(N__30319),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    CascadeMux I__5263 (
            .O(N__30316),
            .I(N__30313));
    InMux I__5262 (
            .O(N__30313),
            .I(N__30308));
    InMux I__5261 (
            .O(N__30312),
            .I(N__30305));
    InMux I__5260 (
            .O(N__30311),
            .I(N__30301));
    LocalMux I__5259 (
            .O(N__30308),
            .I(N__30298));
    LocalMux I__5258 (
            .O(N__30305),
            .I(N__30295));
    InMux I__5257 (
            .O(N__30304),
            .I(N__30292));
    LocalMux I__5256 (
            .O(N__30301),
            .I(N__30288));
    Span4Mux_v I__5255 (
            .O(N__30298),
            .I(N__30281));
    Span4Mux_h I__5254 (
            .O(N__30295),
            .I(N__30281));
    LocalMux I__5253 (
            .O(N__30292),
            .I(N__30281));
    InMux I__5252 (
            .O(N__30291),
            .I(N__30278));
    Span4Mux_v I__5251 (
            .O(N__30288),
            .I(N__30273));
    Span4Mux_h I__5250 (
            .O(N__30281),
            .I(N__30273));
    LocalMux I__5249 (
            .O(N__30278),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__5248 (
            .O(N__30273),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__5247 (
            .O(N__30268),
            .I(N__30265));
    LocalMux I__5246 (
            .O(N__30265),
            .I(\current_shift_inst.control_input_axb_0 ));
    InMux I__5245 (
            .O(N__30262),
            .I(N__30258));
    CascadeMux I__5244 (
            .O(N__30261),
            .I(N__30254));
    LocalMux I__5243 (
            .O(N__30258),
            .I(N__30251));
    InMux I__5242 (
            .O(N__30257),
            .I(N__30248));
    InMux I__5241 (
            .O(N__30254),
            .I(N__30245));
    Span4Mux_h I__5240 (
            .O(N__30251),
            .I(N__30242));
    LocalMux I__5239 (
            .O(N__30248),
            .I(\current_shift_inst.N_1474_i ));
    LocalMux I__5238 (
            .O(N__30245),
            .I(\current_shift_inst.N_1474_i ));
    Odrv4 I__5237 (
            .O(N__30242),
            .I(\current_shift_inst.N_1474_i ));
    InMux I__5236 (
            .O(N__30235),
            .I(N__30232));
    LocalMux I__5235 (
            .O(N__30232),
            .I(N__30229));
    Odrv4 I__5234 (
            .O(N__30229),
            .I(\current_shift_inst.control_input_18 ));
    InMux I__5233 (
            .O(N__30226),
            .I(N__30223));
    LocalMux I__5232 (
            .O(N__30223),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__5231 (
            .O(N__30220),
            .I(N__30217));
    LocalMux I__5230 (
            .O(N__30217),
            .I(N__30214));
    Odrv4 I__5229 (
            .O(N__30214),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__5228 (
            .O(N__30211),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__5227 (
            .O(N__30208),
            .I(N__30205));
    LocalMux I__5226 (
            .O(N__30205),
            .I(N__30202));
    Odrv4 I__5225 (
            .O(N__30202),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__5224 (
            .O(N__30199),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__5223 (
            .O(N__30196),
            .I(N__30193));
    LocalMux I__5222 (
            .O(N__30193),
            .I(N__30190));
    Odrv4 I__5221 (
            .O(N__30190),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__5220 (
            .O(N__30187),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__5219 (
            .O(N__30184),
            .I(N__30181));
    LocalMux I__5218 (
            .O(N__30181),
            .I(N__30178));
    Odrv4 I__5217 (
            .O(N__30178),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__5216 (
            .O(N__30175),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__5215 (
            .O(N__30172),
            .I(N__30169));
    LocalMux I__5214 (
            .O(N__30169),
            .I(N__30166));
    Odrv4 I__5213 (
            .O(N__30166),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__5212 (
            .O(N__30163),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__5211 (
            .O(N__30160),
            .I(N__30157));
    LocalMux I__5210 (
            .O(N__30157),
            .I(N__30154));
    Odrv4 I__5209 (
            .O(N__30154),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__5208 (
            .O(N__30151),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__5207 (
            .O(N__30148),
            .I(N__30143));
    InMux I__5206 (
            .O(N__30147),
            .I(N__30140));
    InMux I__5205 (
            .O(N__30146),
            .I(N__30137));
    LocalMux I__5204 (
            .O(N__30143),
            .I(N__30134));
    LocalMux I__5203 (
            .O(N__30140),
            .I(N__30129));
    LocalMux I__5202 (
            .O(N__30137),
            .I(N__30129));
    Odrv12 I__5201 (
            .O(N__30134),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv12 I__5200 (
            .O(N__30129),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__5199 (
            .O(N__30124),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__5198 (
            .O(N__30121),
            .I(N__30116));
    InMux I__5197 (
            .O(N__30120),
            .I(N__30113));
    InMux I__5196 (
            .O(N__30119),
            .I(N__30110));
    LocalMux I__5195 (
            .O(N__30116),
            .I(N__30105));
    LocalMux I__5194 (
            .O(N__30113),
            .I(N__30105));
    LocalMux I__5193 (
            .O(N__30110),
            .I(N__30102));
    Span4Mux_v I__5192 (
            .O(N__30105),
            .I(N__30099));
    Odrv12 I__5191 (
            .O(N__30102),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv4 I__5190 (
            .O(N__30099),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__5189 (
            .O(N__30094),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    CascadeMux I__5188 (
            .O(N__30091),
            .I(N__30087));
    InMux I__5187 (
            .O(N__30090),
            .I(N__30083));
    InMux I__5186 (
            .O(N__30087),
            .I(N__30080));
    InMux I__5185 (
            .O(N__30086),
            .I(N__30077));
    LocalMux I__5184 (
            .O(N__30083),
            .I(N__30074));
    LocalMux I__5183 (
            .O(N__30080),
            .I(N__30069));
    LocalMux I__5182 (
            .O(N__30077),
            .I(N__30069));
    Odrv4 I__5181 (
            .O(N__30074),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv12 I__5180 (
            .O(N__30069),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__5179 (
            .O(N__30064),
            .I(bfn_12_10_0_));
    InMux I__5178 (
            .O(N__30061),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__5177 (
            .O(N__30058),
            .I(N__30053));
    InMux I__5176 (
            .O(N__30057),
            .I(N__30048));
    InMux I__5175 (
            .O(N__30056),
            .I(N__30048));
    LocalMux I__5174 (
            .O(N__30053),
            .I(N__30045));
    LocalMux I__5173 (
            .O(N__30048),
            .I(N__30042));
    Odrv4 I__5172 (
            .O(N__30045),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv12 I__5171 (
            .O(N__30042),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__5170 (
            .O(N__30037),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__5169 (
            .O(N__30034),
            .I(N__30029));
    InMux I__5168 (
            .O(N__30033),
            .I(N__30024));
    InMux I__5167 (
            .O(N__30032),
            .I(N__30024));
    LocalMux I__5166 (
            .O(N__30029),
            .I(N__30021));
    LocalMux I__5165 (
            .O(N__30024),
            .I(N__30018));
    Odrv4 I__5164 (
            .O(N__30021),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv12 I__5163 (
            .O(N__30018),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__5162 (
            .O(N__30013),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__5161 (
            .O(N__30010),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__5160 (
            .O(N__30007),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__5159 (
            .O(N__30004),
            .I(N__30000));
    InMux I__5158 (
            .O(N__30003),
            .I(N__29994));
    LocalMux I__5157 (
            .O(N__30000),
            .I(N__29991));
    InMux I__5156 (
            .O(N__29999),
            .I(N__29988));
    InMux I__5155 (
            .O(N__29998),
            .I(N__29985));
    InMux I__5154 (
            .O(N__29997),
            .I(N__29982));
    LocalMux I__5153 (
            .O(N__29994),
            .I(N__29979));
    Span4Mux_v I__5152 (
            .O(N__29991),
            .I(N__29974));
    LocalMux I__5151 (
            .O(N__29988),
            .I(N__29974));
    LocalMux I__5150 (
            .O(N__29985),
            .I(N__29971));
    LocalMux I__5149 (
            .O(N__29982),
            .I(N__29968));
    Span4Mux_h I__5148 (
            .O(N__29979),
            .I(N__29963));
    Span4Mux_h I__5147 (
            .O(N__29974),
            .I(N__29963));
    Odrv12 I__5146 (
            .O(N__29971),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__5145 (
            .O(N__29968),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__5144 (
            .O(N__29963),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__5143 (
            .O(N__29956),
            .I(N__29953));
    InMux I__5142 (
            .O(N__29953),
            .I(N__29950));
    LocalMux I__5141 (
            .O(N__29950),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0 ));
    CascadeMux I__5140 (
            .O(N__29947),
            .I(N__29944));
    InMux I__5139 (
            .O(N__29944),
            .I(N__29941));
    LocalMux I__5138 (
            .O(N__29941),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0 ));
    InMux I__5137 (
            .O(N__29938),
            .I(N__29935));
    LocalMux I__5136 (
            .O(N__29935),
            .I(\current_shift_inst.PI_CTRL.integrator_i_20 ));
    InMux I__5135 (
            .O(N__29932),
            .I(N__29929));
    LocalMux I__5134 (
            .O(N__29929),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__5133 (
            .O(N__29926),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__5132 (
            .O(N__29923),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__5131 (
            .O(N__29920),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    CascadeMux I__5130 (
            .O(N__29917),
            .I(N__29913));
    InMux I__5129 (
            .O(N__29916),
            .I(N__29909));
    InMux I__5128 (
            .O(N__29913),
            .I(N__29906));
    InMux I__5127 (
            .O(N__29912),
            .I(N__29903));
    LocalMux I__5126 (
            .O(N__29909),
            .I(N__29900));
    LocalMux I__5125 (
            .O(N__29906),
            .I(N__29895));
    LocalMux I__5124 (
            .O(N__29903),
            .I(N__29895));
    Odrv12 I__5123 (
            .O(N__29900),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv12 I__5122 (
            .O(N__29895),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__5121 (
            .O(N__29890),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    CascadeMux I__5120 (
            .O(N__29887),
            .I(N__29883));
    InMux I__5119 (
            .O(N__29886),
            .I(N__29879));
    InMux I__5118 (
            .O(N__29883),
            .I(N__29876));
    InMux I__5117 (
            .O(N__29882),
            .I(N__29873));
    LocalMux I__5116 (
            .O(N__29879),
            .I(N__29870));
    LocalMux I__5115 (
            .O(N__29876),
            .I(N__29865));
    LocalMux I__5114 (
            .O(N__29873),
            .I(N__29865));
    Odrv12 I__5113 (
            .O(N__29870),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv12 I__5112 (
            .O(N__29865),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__5111 (
            .O(N__29860),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    CascadeMux I__5110 (
            .O(N__29857),
            .I(N__29853));
    InMux I__5109 (
            .O(N__29856),
            .I(N__29849));
    InMux I__5108 (
            .O(N__29853),
            .I(N__29846));
    CascadeMux I__5107 (
            .O(N__29852),
            .I(N__29843));
    LocalMux I__5106 (
            .O(N__29849),
            .I(N__29838));
    LocalMux I__5105 (
            .O(N__29846),
            .I(N__29835));
    InMux I__5104 (
            .O(N__29843),
            .I(N__29832));
    CascadeMux I__5103 (
            .O(N__29842),
            .I(N__29829));
    InMux I__5102 (
            .O(N__29841),
            .I(N__29826));
    Span4Mux_h I__5101 (
            .O(N__29838),
            .I(N__29821));
    Span4Mux_h I__5100 (
            .O(N__29835),
            .I(N__29821));
    LocalMux I__5099 (
            .O(N__29832),
            .I(N__29818));
    InMux I__5098 (
            .O(N__29829),
            .I(N__29815));
    LocalMux I__5097 (
            .O(N__29826),
            .I(N__29812));
    Odrv4 I__5096 (
            .O(N__29821),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv12 I__5095 (
            .O(N__29818),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__5094 (
            .O(N__29815),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__5093 (
            .O(N__29812),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__5092 (
            .O(N__29803),
            .I(N__29800));
    LocalMux I__5091 (
            .O(N__29800),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0 ));
    CascadeMux I__5090 (
            .O(N__29797),
            .I(N__29794));
    InMux I__5089 (
            .O(N__29794),
            .I(N__29790));
    InMux I__5088 (
            .O(N__29793),
            .I(N__29786));
    LocalMux I__5087 (
            .O(N__29790),
            .I(N__29781));
    InMux I__5086 (
            .O(N__29789),
            .I(N__29778));
    LocalMux I__5085 (
            .O(N__29786),
            .I(N__29775));
    InMux I__5084 (
            .O(N__29785),
            .I(N__29770));
    InMux I__5083 (
            .O(N__29784),
            .I(N__29770));
    Span4Mux_h I__5082 (
            .O(N__29781),
            .I(N__29767));
    LocalMux I__5081 (
            .O(N__29778),
            .I(N__29760));
    Span4Mux_h I__5080 (
            .O(N__29775),
            .I(N__29760));
    LocalMux I__5079 (
            .O(N__29770),
            .I(N__29760));
    Odrv4 I__5078 (
            .O(N__29767),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__5077 (
            .O(N__29760),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__5076 (
            .O(N__29755),
            .I(N__29752));
    InMux I__5075 (
            .O(N__29752),
            .I(N__29749));
    LocalMux I__5074 (
            .O(N__29749),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0 ));
    CascadeMux I__5073 (
            .O(N__29746),
            .I(N__29743));
    InMux I__5072 (
            .O(N__29743),
            .I(N__29740));
    LocalMux I__5071 (
            .O(N__29740),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0 ));
    CascadeMux I__5070 (
            .O(N__29737),
            .I(N__29734));
    InMux I__5069 (
            .O(N__29734),
            .I(N__29731));
    LocalMux I__5068 (
            .O(N__29731),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0 ));
    CascadeMux I__5067 (
            .O(N__29728),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25_cascade_ ));
    InMux I__5066 (
            .O(N__29725),
            .I(N__29722));
    LocalMux I__5065 (
            .O(N__29722),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0 ));
    InMux I__5064 (
            .O(N__29719),
            .I(N__29715));
    InMux I__5063 (
            .O(N__29718),
            .I(N__29711));
    LocalMux I__5062 (
            .O(N__29715),
            .I(N__29708));
    InMux I__5061 (
            .O(N__29714),
            .I(N__29705));
    LocalMux I__5060 (
            .O(N__29711),
            .I(N__29700));
    Span4Mux_h I__5059 (
            .O(N__29708),
            .I(N__29695));
    LocalMux I__5058 (
            .O(N__29705),
            .I(N__29695));
    InMux I__5057 (
            .O(N__29704),
            .I(N__29692));
    InMux I__5056 (
            .O(N__29703),
            .I(N__29689));
    Span4Mux_h I__5055 (
            .O(N__29700),
            .I(N__29682));
    Span4Mux_h I__5054 (
            .O(N__29695),
            .I(N__29682));
    LocalMux I__5053 (
            .O(N__29692),
            .I(N__29682));
    LocalMux I__5052 (
            .O(N__29689),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__5051 (
            .O(N__29682),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    CascadeMux I__5050 (
            .O(N__29677),
            .I(N__29674));
    InMux I__5049 (
            .O(N__29674),
            .I(N__29671));
    LocalMux I__5048 (
            .O(N__29671),
            .I(N__29668));
    Odrv4 I__5047 (
            .O(N__29668),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0 ));
    CascadeMux I__5046 (
            .O(N__29665),
            .I(N__29662));
    InMux I__5045 (
            .O(N__29662),
            .I(N__29659));
    LocalMux I__5044 (
            .O(N__29659),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0 ));
    CascadeMux I__5043 (
            .O(N__29656),
            .I(N__29653));
    InMux I__5042 (
            .O(N__29653),
            .I(N__29649));
    InMux I__5041 (
            .O(N__29652),
            .I(N__29646));
    LocalMux I__5040 (
            .O(N__29649),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_14 ));
    LocalMux I__5039 (
            .O(N__29646),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_14 ));
    CascadeMux I__5038 (
            .O(N__29641),
            .I(N__29638));
    InMux I__5037 (
            .O(N__29638),
            .I(N__29634));
    InMux I__5036 (
            .O(N__29637),
            .I(N__29630));
    LocalMux I__5035 (
            .O(N__29634),
            .I(N__29627));
    InMux I__5034 (
            .O(N__29633),
            .I(N__29624));
    LocalMux I__5033 (
            .O(N__29630),
            .I(N__29620));
    Span4Mux_v I__5032 (
            .O(N__29627),
            .I(N__29615));
    LocalMux I__5031 (
            .O(N__29624),
            .I(N__29615));
    InMux I__5030 (
            .O(N__29623),
            .I(N__29611));
    Span4Mux_h I__5029 (
            .O(N__29620),
            .I(N__29608));
    Span4Mux_h I__5028 (
            .O(N__29615),
            .I(N__29605));
    InMux I__5027 (
            .O(N__29614),
            .I(N__29602));
    LocalMux I__5026 (
            .O(N__29611),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__5025 (
            .O(N__29608),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__5024 (
            .O(N__29605),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__5023 (
            .O(N__29602),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__5022 (
            .O(N__29593),
            .I(N__29590));
    LocalMux I__5021 (
            .O(N__29590),
            .I(\current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9 ));
    CascadeMux I__5020 (
            .O(N__29587),
            .I(N__29584));
    InMux I__5019 (
            .O(N__29584),
            .I(N__29579));
    InMux I__5018 (
            .O(N__29583),
            .I(N__29576));
    InMux I__5017 (
            .O(N__29582),
            .I(N__29573));
    LocalMux I__5016 (
            .O(N__29579),
            .I(N__29570));
    LocalMux I__5015 (
            .O(N__29576),
            .I(N__29567));
    LocalMux I__5014 (
            .O(N__29573),
            .I(N__29563));
    Span4Mux_v I__5013 (
            .O(N__29570),
            .I(N__29560));
    Span4Mux_h I__5012 (
            .O(N__29567),
            .I(N__29556));
    InMux I__5011 (
            .O(N__29566),
            .I(N__29553));
    Span4Mux_h I__5010 (
            .O(N__29563),
            .I(N__29550));
    Span4Mux_h I__5009 (
            .O(N__29560),
            .I(N__29547));
    InMux I__5008 (
            .O(N__29559),
            .I(N__29544));
    Odrv4 I__5007 (
            .O(N__29556),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__5006 (
            .O(N__29553),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__5005 (
            .O(N__29550),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__5004 (
            .O(N__29547),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__5003 (
            .O(N__29544),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__5002 (
            .O(N__29533),
            .I(N__29530));
    InMux I__5001 (
            .O(N__29530),
            .I(N__29527));
    LocalMux I__5000 (
            .O(N__29527),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8 ));
    CascadeMux I__4999 (
            .O(N__29524),
            .I(N__29521));
    InMux I__4998 (
            .O(N__29521),
            .I(N__29518));
    LocalMux I__4997 (
            .O(N__29518),
            .I(N__29515));
    Odrv4 I__4996 (
            .O(N__29515),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0 ));
    CascadeMux I__4995 (
            .O(N__29512),
            .I(N__29509));
    InMux I__4994 (
            .O(N__29509),
            .I(N__29506));
    LocalMux I__4993 (
            .O(N__29506),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0 ));
    InMux I__4992 (
            .O(N__29503),
            .I(N__29500));
    LocalMux I__4991 (
            .O(N__29500),
            .I(\current_shift_inst.PI_CTRL.integrator_i_10 ));
    InMux I__4990 (
            .O(N__29497),
            .I(N__29494));
    LocalMux I__4989 (
            .O(N__29494),
            .I(\current_shift_inst.PI_CTRL.integrator_i_13 ));
    InMux I__4988 (
            .O(N__29491),
            .I(N__29487));
    InMux I__4987 (
            .O(N__29490),
            .I(N__29484));
    LocalMux I__4986 (
            .O(N__29487),
            .I(N__29478));
    LocalMux I__4985 (
            .O(N__29484),
            .I(N__29475));
    CascadeMux I__4984 (
            .O(N__29483),
            .I(N__29472));
    CascadeMux I__4983 (
            .O(N__29482),
            .I(N__29469));
    InMux I__4982 (
            .O(N__29481),
            .I(N__29466));
    Span4Mux_h I__4981 (
            .O(N__29478),
            .I(N__29463));
    Span4Mux_h I__4980 (
            .O(N__29475),
            .I(N__29460));
    InMux I__4979 (
            .O(N__29472),
            .I(N__29455));
    InMux I__4978 (
            .O(N__29469),
            .I(N__29455));
    LocalMux I__4977 (
            .O(N__29466),
            .I(N__29452));
    Odrv4 I__4976 (
            .O(N__29463),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__4975 (
            .O(N__29460),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__4974 (
            .O(N__29455),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__4973 (
            .O(N__29452),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__4972 (
            .O(N__29443),
            .I(N__29440));
    InMux I__4971 (
            .O(N__29440),
            .I(N__29437));
    LocalMux I__4970 (
            .O(N__29437),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0 ));
    CascadeMux I__4969 (
            .O(N__29434),
            .I(N__29431));
    InMux I__4968 (
            .O(N__29431),
            .I(N__29427));
    InMux I__4967 (
            .O(N__29430),
            .I(N__29424));
    LocalMux I__4966 (
            .O(N__29427),
            .I(N__29421));
    LocalMux I__4965 (
            .O(N__29424),
            .I(N__29417));
    Span4Mux_v I__4964 (
            .O(N__29421),
            .I(N__29413));
    InMux I__4963 (
            .O(N__29420),
            .I(N__29410));
    Span4Mux_v I__4962 (
            .O(N__29417),
            .I(N__29407));
    InMux I__4961 (
            .O(N__29416),
            .I(N__29404));
    Span4Mux_h I__4960 (
            .O(N__29413),
            .I(N__29401));
    LocalMux I__4959 (
            .O(N__29410),
            .I(N__29398));
    Odrv4 I__4958 (
            .O(N__29407),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__4957 (
            .O(N__29404),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__4956 (
            .O(N__29401),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__4955 (
            .O(N__29398),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__4954 (
            .O(N__29389),
            .I(N__29386));
    InMux I__4953 (
            .O(N__29386),
            .I(N__29383));
    LocalMux I__4952 (
            .O(N__29383),
            .I(N__29380));
    Odrv4 I__4951 (
            .O(N__29380),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5 ));
    InMux I__4950 (
            .O(N__29377),
            .I(N__29374));
    LocalMux I__4949 (
            .O(N__29374),
            .I(N__29370));
    InMux I__4948 (
            .O(N__29373),
            .I(N__29367));
    Span4Mux_v I__4947 (
            .O(N__29370),
            .I(N__29364));
    LocalMux I__4946 (
            .O(N__29367),
            .I(N__29361));
    Odrv4 I__4945 (
            .O(N__29364),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    Odrv12 I__4944 (
            .O(N__29361),
            .I(\current_shift_inst.PI_CTRL.integrator_i_0 ));
    CascadeMux I__4943 (
            .O(N__29356),
            .I(N__29353));
    InMux I__4942 (
            .O(N__29353),
            .I(N__29350));
    LocalMux I__4941 (
            .O(N__29350),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4 ));
    CascadeMux I__4940 (
            .O(N__29347),
            .I(N__29343));
    CascadeMux I__4939 (
            .O(N__29346),
            .I(N__29340));
    InMux I__4938 (
            .O(N__29343),
            .I(N__29335));
    InMux I__4937 (
            .O(N__29340),
            .I(N__29332));
    InMux I__4936 (
            .O(N__29339),
            .I(N__29329));
    InMux I__4935 (
            .O(N__29338),
            .I(N__29325));
    LocalMux I__4934 (
            .O(N__29335),
            .I(N__29322));
    LocalMux I__4933 (
            .O(N__29332),
            .I(N__29319));
    LocalMux I__4932 (
            .O(N__29329),
            .I(N__29316));
    InMux I__4931 (
            .O(N__29328),
            .I(N__29313));
    LocalMux I__4930 (
            .O(N__29325),
            .I(N__29310));
    Span4Mux_h I__4929 (
            .O(N__29322),
            .I(N__29307));
    Span4Mux_h I__4928 (
            .O(N__29319),
            .I(N__29304));
    Span4Mux_h I__4927 (
            .O(N__29316),
            .I(N__29297));
    LocalMux I__4926 (
            .O(N__29313),
            .I(N__29297));
    Span4Mux_h I__4925 (
            .O(N__29310),
            .I(N__29297));
    Odrv4 I__4924 (
            .O(N__29307),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__4923 (
            .O(N__29304),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__4922 (
            .O(N__29297),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__4921 (
            .O(N__29290),
            .I(N__29287));
    InMux I__4920 (
            .O(N__29287),
            .I(N__29284));
    LocalMux I__4919 (
            .O(N__29284),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10 ));
    CascadeMux I__4918 (
            .O(N__29281),
            .I(N__29278));
    InMux I__4917 (
            .O(N__29278),
            .I(N__29275));
    LocalMux I__4916 (
            .O(N__29275),
            .I(N__29272));
    Span4Mux_h I__4915 (
            .O(N__29272),
            .I(N__29269));
    Odrv4 I__4914 (
            .O(N__29269),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13 ));
    InMux I__4913 (
            .O(N__29266),
            .I(N__29263));
    LocalMux I__4912 (
            .O(N__29263),
            .I(N__29258));
    InMux I__4911 (
            .O(N__29262),
            .I(N__29254));
    InMux I__4910 (
            .O(N__29261),
            .I(N__29251));
    Span4Mux_h I__4909 (
            .O(N__29258),
            .I(N__29248));
    InMux I__4908 (
            .O(N__29257),
            .I(N__29245));
    LocalMux I__4907 (
            .O(N__29254),
            .I(N__29242));
    LocalMux I__4906 (
            .O(N__29251),
            .I(N__29239));
    Span4Mux_h I__4905 (
            .O(N__29248),
            .I(N__29234));
    LocalMux I__4904 (
            .O(N__29245),
            .I(N__29234));
    Span4Mux_v I__4903 (
            .O(N__29242),
            .I(N__29229));
    Span4Mux_h I__4902 (
            .O(N__29239),
            .I(N__29229));
    Odrv4 I__4901 (
            .O(N__29234),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__4900 (
            .O(N__29229),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    CascadeMux I__4899 (
            .O(N__29224),
            .I(N__29221));
    InMux I__4898 (
            .O(N__29221),
            .I(N__29218));
    LocalMux I__4897 (
            .O(N__29218),
            .I(\current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6 ));
    CascadeMux I__4896 (
            .O(N__29215),
            .I(N__29211));
    InMux I__4895 (
            .O(N__29214),
            .I(N__29208));
    InMux I__4894 (
            .O(N__29211),
            .I(N__29205));
    LocalMux I__4893 (
            .O(N__29208),
            .I(N__29200));
    LocalMux I__4892 (
            .O(N__29205),
            .I(N__29197));
    InMux I__4891 (
            .O(N__29204),
            .I(N__29194));
    InMux I__4890 (
            .O(N__29203),
            .I(N__29190));
    Span4Mux_v I__4889 (
            .O(N__29200),
            .I(N__29183));
    Span4Mux_v I__4888 (
            .O(N__29197),
            .I(N__29183));
    LocalMux I__4887 (
            .O(N__29194),
            .I(N__29183));
    InMux I__4886 (
            .O(N__29193),
            .I(N__29180));
    LocalMux I__4885 (
            .O(N__29190),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__4884 (
            .O(N__29183),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__4883 (
            .O(N__29180),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    CascadeMux I__4882 (
            .O(N__29173),
            .I(N__29170));
    InMux I__4881 (
            .O(N__29170),
            .I(N__29167));
    LocalMux I__4880 (
            .O(N__29167),
            .I(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0 ));
    CascadeMux I__4879 (
            .O(N__29164),
            .I(N__29161));
    InMux I__4878 (
            .O(N__29161),
            .I(N__29158));
    LocalMux I__4877 (
            .O(N__29158),
            .I(\current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11 ));
    InMux I__4876 (
            .O(N__29155),
            .I(N__29151));
    InMux I__4875 (
            .O(N__29154),
            .I(N__29148));
    LocalMux I__4874 (
            .O(N__29151),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__4873 (
            .O(N__29148),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__4872 (
            .O(N__29143),
            .I(N__29139));
    InMux I__4871 (
            .O(N__29142),
            .I(N__29136));
    LocalMux I__4870 (
            .O(N__29139),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__4869 (
            .O(N__29136),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__4868 (
            .O(N__29131),
            .I(N__29128));
    LocalMux I__4867 (
            .O(N__29128),
            .I(N__29125));
    Odrv12 I__4866 (
            .O(N__29125),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df28 ));
    CascadeMux I__4865 (
            .O(N__29122),
            .I(N__29119));
    InMux I__4864 (
            .O(N__29119),
            .I(N__29116));
    LocalMux I__4863 (
            .O(N__29116),
            .I(N__29110));
    InMux I__4862 (
            .O(N__29115),
            .I(N__29107));
    InMux I__4861 (
            .O(N__29114),
            .I(N__29104));
    InMux I__4860 (
            .O(N__29113),
            .I(N__29101));
    Span4Mux_h I__4859 (
            .O(N__29110),
            .I(N__29096));
    LocalMux I__4858 (
            .O(N__29107),
            .I(N__29096));
    LocalMux I__4857 (
            .O(N__29104),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    LocalMux I__4856 (
            .O(N__29101),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv4 I__4855 (
            .O(N__29096),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__4854 (
            .O(N__29089),
            .I(N__29084));
    InMux I__4853 (
            .O(N__29088),
            .I(N__29081));
    InMux I__4852 (
            .O(N__29087),
            .I(N__29078));
    LocalMux I__4851 (
            .O(N__29084),
            .I(N__29075));
    LocalMux I__4850 (
            .O(N__29081),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__4849 (
            .O(N__29078),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__4848 (
            .O(N__29075),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__4847 (
            .O(N__29068),
            .I(N__29065));
    LocalMux I__4846 (
            .O(N__29065),
            .I(N__29062));
    Odrv4 I__4845 (
            .O(N__29062),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    InMux I__4844 (
            .O(N__29059),
            .I(N__29056));
    LocalMux I__4843 (
            .O(N__29056),
            .I(N__29052));
    InMux I__4842 (
            .O(N__29055),
            .I(N__29049));
    Span12Mux_v I__4841 (
            .O(N__29052),
            .I(N__29044));
    LocalMux I__4840 (
            .O(N__29049),
            .I(N__29041));
    InMux I__4839 (
            .O(N__29048),
            .I(N__29038));
    InMux I__4838 (
            .O(N__29047),
            .I(N__29035));
    Span12Mux_v I__4837 (
            .O(N__29044),
            .I(N__29032));
    Span12Mux_v I__4836 (
            .O(N__29041),
            .I(N__29029));
    LocalMux I__4835 (
            .O(N__29038),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__4834 (
            .O(N__29035),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv12 I__4833 (
            .O(N__29032),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv12 I__4832 (
            .O(N__29029),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__4831 (
            .O(N__29020),
            .I(N__29014));
    ClkMux I__4830 (
            .O(N__29019),
            .I(N__29014));
    GlobalMux I__4829 (
            .O(N__29014),
            .I(N__29011));
    gio2CtrlBuf I__4828 (
            .O(N__29011),
            .I(delay_tr_input_c_g));
    InMux I__4827 (
            .O(N__29008),
            .I(N__29005));
    LocalMux I__4826 (
            .O(N__29005),
            .I(N__29002));
    Span4Mux_v I__4825 (
            .O(N__29002),
            .I(N__28999));
    Span4Mux_v I__4824 (
            .O(N__28999),
            .I(N__28994));
    InMux I__4823 (
            .O(N__28998),
            .I(N__28991));
    InMux I__4822 (
            .O(N__28997),
            .I(N__28988));
    Span4Mux_v I__4821 (
            .O(N__28994),
            .I(N__28985));
    LocalMux I__4820 (
            .O(N__28991),
            .I(N__28982));
    LocalMux I__4819 (
            .O(N__28988),
            .I(N__28979));
    Span4Mux_v I__4818 (
            .O(N__28985),
            .I(N__28976));
    Sp12to4 I__4817 (
            .O(N__28982),
            .I(N__28973));
    Span12Mux_v I__4816 (
            .O(N__28979),
            .I(N__28970));
    Span4Mux_v I__4815 (
            .O(N__28976),
            .I(N__28967));
    Odrv12 I__4814 (
            .O(N__28973),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv12 I__4813 (
            .O(N__28970),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    Odrv4 I__4812 (
            .O(N__28967),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    IoInMux I__4811 (
            .O(N__28960),
            .I(N__28957));
    LocalMux I__4810 (
            .O(N__28957),
            .I(N__28954));
    Odrv4 I__4809 (
            .O(N__28954),
            .I(\delay_measurement_inst.delay_tr_timer.N_399_i ));
    CascadeMux I__4808 (
            .O(N__28951),
            .I(N__28948));
    InMux I__4807 (
            .O(N__28948),
            .I(N__28945));
    LocalMux I__4806 (
            .O(N__28945),
            .I(N__28942));
    Odrv4 I__4805 (
            .O(N__28942),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__4804 (
            .O(N__28939),
            .I(N__28933));
    InMux I__4803 (
            .O(N__28938),
            .I(N__28933));
    LocalMux I__4802 (
            .O(N__28933),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__4801 (
            .O(N__28930),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    InMux I__4800 (
            .O(N__28927),
            .I(N__28924));
    LocalMux I__4799 (
            .O(N__28924),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    InMux I__4798 (
            .O(N__28921),
            .I(N__28909));
    InMux I__4797 (
            .O(N__28920),
            .I(N__28909));
    InMux I__4796 (
            .O(N__28919),
            .I(N__28909));
    InMux I__4795 (
            .O(N__28918),
            .I(N__28909));
    LocalMux I__4794 (
            .O(N__28909),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__4793 (
            .O(N__28906),
            .I(N__28902));
    CascadeMux I__4792 (
            .O(N__28905),
            .I(N__28899));
    InMux I__4791 (
            .O(N__28902),
            .I(N__28894));
    InMux I__4790 (
            .O(N__28899),
            .I(N__28894));
    LocalMux I__4789 (
            .O(N__28894),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__4788 (
            .O(N__28891),
            .I(N__28888));
    LocalMux I__4787 (
            .O(N__28888),
            .I(N__28885));
    Odrv4 I__4786 (
            .O(N__28885),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    InMux I__4785 (
            .O(N__28882),
            .I(N__28878));
    InMux I__4784 (
            .O(N__28881),
            .I(N__28875));
    LocalMux I__4783 (
            .O(N__28878),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    LocalMux I__4782 (
            .O(N__28875),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__4781 (
            .O(N__28870),
            .I(N__28866));
    InMux I__4780 (
            .O(N__28869),
            .I(N__28863));
    LocalMux I__4779 (
            .O(N__28866),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    LocalMux I__4778 (
            .O(N__28863),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__4777 (
            .O(N__28858),
            .I(N__28855));
    LocalMux I__4776 (
            .O(N__28855),
            .I(N__28852));
    Odrv4 I__4775 (
            .O(N__28852),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df20 ));
    InMux I__4774 (
            .O(N__28849),
            .I(N__28845));
    InMux I__4773 (
            .O(N__28848),
            .I(N__28842));
    LocalMux I__4772 (
            .O(N__28845),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    LocalMux I__4771 (
            .O(N__28842),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__4770 (
            .O(N__28837),
            .I(N__28833));
    InMux I__4769 (
            .O(N__28836),
            .I(N__28830));
    LocalMux I__4768 (
            .O(N__28833),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    LocalMux I__4767 (
            .O(N__28830),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__4766 (
            .O(N__28825),
            .I(N__28822));
    LocalMux I__4765 (
            .O(N__28822),
            .I(N__28819));
    Odrv4 I__4764 (
            .O(N__28819),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df22 ));
    InMux I__4763 (
            .O(N__28816),
            .I(N__28812));
    InMux I__4762 (
            .O(N__28815),
            .I(N__28809));
    LocalMux I__4761 (
            .O(N__28812),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__4760 (
            .O(N__28809),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__4759 (
            .O(N__28804),
            .I(N__28800));
    InMux I__4758 (
            .O(N__28803),
            .I(N__28797));
    LocalMux I__4757 (
            .O(N__28800),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__4756 (
            .O(N__28797),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__4755 (
            .O(N__28792),
            .I(N__28789));
    LocalMux I__4754 (
            .O(N__28789),
            .I(N__28786));
    Odrv4 I__4753 (
            .O(N__28786),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df24 ));
    InMux I__4752 (
            .O(N__28783),
            .I(N__28779));
    InMux I__4751 (
            .O(N__28782),
            .I(N__28776));
    LocalMux I__4750 (
            .O(N__28779),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__4749 (
            .O(N__28776),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__4748 (
            .O(N__28771),
            .I(N__28767));
    InMux I__4747 (
            .O(N__28770),
            .I(N__28764));
    LocalMux I__4746 (
            .O(N__28767),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__4745 (
            .O(N__28764),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__4744 (
            .O(N__28759),
            .I(N__28756));
    LocalMux I__4743 (
            .O(N__28756),
            .I(N__28753));
    Odrv4 I__4742 (
            .O(N__28753),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df26 ));
    InMux I__4741 (
            .O(N__28750),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ));
    InMux I__4740 (
            .O(N__28747),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    CascadeMux I__4739 (
            .O(N__28744),
            .I(N__28741));
    InMux I__4738 (
            .O(N__28741),
            .I(N__28738));
    LocalMux I__4737 (
            .O(N__28738),
            .I(N__28735));
    Odrv4 I__4736 (
            .O(N__28735),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28 ));
    InMux I__4735 (
            .O(N__28732),
            .I(N__28726));
    InMux I__4734 (
            .O(N__28731),
            .I(N__28726));
    LocalMux I__4733 (
            .O(N__28726),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    CascadeMux I__4732 (
            .O(N__28723),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ));
    CascadeMux I__4731 (
            .O(N__28720),
            .I(N__28715));
    InMux I__4730 (
            .O(N__28719),
            .I(N__28712));
    InMux I__4729 (
            .O(N__28718),
            .I(N__28709));
    InMux I__4728 (
            .O(N__28715),
            .I(N__28706));
    LocalMux I__4727 (
            .O(N__28712),
            .I(N__28703));
    LocalMux I__4726 (
            .O(N__28709),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__4725 (
            .O(N__28706),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__4724 (
            .O(N__28703),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__4723 (
            .O(N__28696),
            .I(N__28692));
    InMux I__4722 (
            .O(N__28695),
            .I(N__28689));
    LocalMux I__4721 (
            .O(N__28692),
            .I(N__28686));
    LocalMux I__4720 (
            .O(N__28689),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__4719 (
            .O(N__28686),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__4718 (
            .O(N__28681),
            .I(N__28678));
    InMux I__4717 (
            .O(N__28678),
            .I(N__28675));
    LocalMux I__4716 (
            .O(N__28675),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__4715 (
            .O(N__28672),
            .I(N__28668));
    InMux I__4714 (
            .O(N__28671),
            .I(N__28665));
    LocalMux I__4713 (
            .O(N__28668),
            .I(N__28662));
    LocalMux I__4712 (
            .O(N__28665),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__4711 (
            .O(N__28662),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__4710 (
            .O(N__28657),
            .I(N__28654));
    InMux I__4709 (
            .O(N__28654),
            .I(N__28651));
    LocalMux I__4708 (
            .O(N__28651),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__4707 (
            .O(N__28648),
            .I(N__28644));
    InMux I__4706 (
            .O(N__28647),
            .I(N__28641));
    LocalMux I__4705 (
            .O(N__28644),
            .I(N__28638));
    LocalMux I__4704 (
            .O(N__28641),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__4703 (
            .O(N__28638),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__4702 (
            .O(N__28633),
            .I(N__28630));
    InMux I__4701 (
            .O(N__28630),
            .I(N__28627));
    LocalMux I__4700 (
            .O(N__28627),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__4699 (
            .O(N__28624),
            .I(N__28620));
    InMux I__4698 (
            .O(N__28623),
            .I(N__28617));
    LocalMux I__4697 (
            .O(N__28620),
            .I(N__28614));
    LocalMux I__4696 (
            .O(N__28617),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__4695 (
            .O(N__28614),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__4694 (
            .O(N__28609),
            .I(N__28606));
    InMux I__4693 (
            .O(N__28606),
            .I(N__28603));
    LocalMux I__4692 (
            .O(N__28603),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__4691 (
            .O(N__28600),
            .I(N__28596));
    InMux I__4690 (
            .O(N__28599),
            .I(N__28593));
    LocalMux I__4689 (
            .O(N__28596),
            .I(N__28590));
    LocalMux I__4688 (
            .O(N__28593),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__4687 (
            .O(N__28590),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__4686 (
            .O(N__28585),
            .I(N__28582));
    LocalMux I__4685 (
            .O(N__28582),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__4684 (
            .O(N__28579),
            .I(N__28575));
    InMux I__4683 (
            .O(N__28578),
            .I(N__28572));
    LocalMux I__4682 (
            .O(N__28575),
            .I(N__28569));
    LocalMux I__4681 (
            .O(N__28572),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__4680 (
            .O(N__28569),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__4679 (
            .O(N__28564),
            .I(N__28561));
    InMux I__4678 (
            .O(N__28561),
            .I(N__28558));
    LocalMux I__4677 (
            .O(N__28558),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__4676 (
            .O(N__28555),
            .I(N__28551));
    InMux I__4675 (
            .O(N__28554),
            .I(N__28548));
    LocalMux I__4674 (
            .O(N__28551),
            .I(N__28545));
    LocalMux I__4673 (
            .O(N__28548),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__4672 (
            .O(N__28545),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__4671 (
            .O(N__28540),
            .I(N__28537));
    LocalMux I__4670 (
            .O(N__28537),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__4669 (
            .O(N__28534),
            .I(N__28530));
    InMux I__4668 (
            .O(N__28533),
            .I(N__28527));
    LocalMux I__4667 (
            .O(N__28530),
            .I(N__28524));
    LocalMux I__4666 (
            .O(N__28527),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__4665 (
            .O(N__28524),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__4664 (
            .O(N__28519),
            .I(N__28516));
    InMux I__4663 (
            .O(N__28516),
            .I(N__28513));
    LocalMux I__4662 (
            .O(N__28513),
            .I(N__28510));
    Odrv4 I__4661 (
            .O(N__28510),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__4660 (
            .O(N__28507),
            .I(N__28503));
    InMux I__4659 (
            .O(N__28506),
            .I(N__28500));
    LocalMux I__4658 (
            .O(N__28503),
            .I(N__28497));
    LocalMux I__4657 (
            .O(N__28500),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__4656 (
            .O(N__28497),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__4655 (
            .O(N__28492),
            .I(N__28489));
    InMux I__4654 (
            .O(N__28489),
            .I(N__28486));
    LocalMux I__4653 (
            .O(N__28486),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__4652 (
            .O(N__28483),
            .I(N__28479));
    InMux I__4651 (
            .O(N__28482),
            .I(N__28476));
    LocalMux I__4650 (
            .O(N__28479),
            .I(N__28473));
    LocalMux I__4649 (
            .O(N__28476),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__4648 (
            .O(N__28473),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__4647 (
            .O(N__28468),
            .I(N__28465));
    LocalMux I__4646 (
            .O(N__28465),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__4645 (
            .O(N__28462),
            .I(N__28458));
    InMux I__4644 (
            .O(N__28461),
            .I(N__28455));
    LocalMux I__4643 (
            .O(N__28458),
            .I(N__28452));
    LocalMux I__4642 (
            .O(N__28455),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__4641 (
            .O(N__28452),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__4640 (
            .O(N__28447),
            .I(N__28444));
    InMux I__4639 (
            .O(N__28444),
            .I(N__28441));
    LocalMux I__4638 (
            .O(N__28441),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__4637 (
            .O(N__28438),
            .I(N__28435));
    LocalMux I__4636 (
            .O(N__28435),
            .I(N__28431));
    InMux I__4635 (
            .O(N__28434),
            .I(N__28428));
    Span4Mux_h I__4634 (
            .O(N__28431),
            .I(N__28425));
    LocalMux I__4633 (
            .O(N__28428),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__4632 (
            .O(N__28425),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__4631 (
            .O(N__28420),
            .I(N__28417));
    InMux I__4630 (
            .O(N__28417),
            .I(N__28414));
    LocalMux I__4629 (
            .O(N__28414),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__4628 (
            .O(N__28411),
            .I(N__28407));
    InMux I__4627 (
            .O(N__28410),
            .I(N__28404));
    LocalMux I__4626 (
            .O(N__28407),
            .I(N__28401));
    LocalMux I__4625 (
            .O(N__28404),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__4624 (
            .O(N__28401),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__4623 (
            .O(N__28396),
            .I(N__28393));
    InMux I__4622 (
            .O(N__28393),
            .I(N__28390));
    LocalMux I__4621 (
            .O(N__28390),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__4620 (
            .O(N__28387),
            .I(N__28384));
    InMux I__4619 (
            .O(N__28384),
            .I(N__28381));
    LocalMux I__4618 (
            .O(N__28381),
            .I(N__28378));
    Span4Mux_h I__4617 (
            .O(N__28378),
            .I(N__28375));
    Odrv4 I__4616 (
            .O(N__28375),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__4615 (
            .O(N__28372),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__4614 (
            .O(N__28369),
            .I(N__28366));
    LocalMux I__4613 (
            .O(N__28366),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__4612 (
            .O(N__28363),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    CascadeMux I__4611 (
            .O(N__28360),
            .I(N__28357));
    InMux I__4610 (
            .O(N__28357),
            .I(N__28354));
    LocalMux I__4609 (
            .O(N__28354),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__4608 (
            .O(N__28351),
            .I(N__28348));
    LocalMux I__4607 (
            .O(N__28348),
            .I(N__28345));
    Odrv12 I__4606 (
            .O(N__28345),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__4605 (
            .O(N__28342),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__4604 (
            .O(N__28339),
            .I(N__28336));
    LocalMux I__4603 (
            .O(N__28336),
            .I(N__28333));
    Span4Mux_v I__4602 (
            .O(N__28333),
            .I(N__28330));
    Odrv4 I__4601 (
            .O(N__28330),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__4600 (
            .O(N__28327),
            .I(N__28324));
    LocalMux I__4599 (
            .O(N__28324),
            .I(N__28321));
    Odrv4 I__4598 (
            .O(N__28321),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__4597 (
            .O(N__28318),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__4596 (
            .O(N__28315),
            .I(N__28305));
    InMux I__4595 (
            .O(N__28314),
            .I(N__28297));
    InMux I__4594 (
            .O(N__28313),
            .I(N__28290));
    InMux I__4593 (
            .O(N__28312),
            .I(N__28290));
    InMux I__4592 (
            .O(N__28311),
            .I(N__28290));
    CascadeMux I__4591 (
            .O(N__28310),
            .I(N__28278));
    InMux I__4590 (
            .O(N__28309),
            .I(N__28263));
    InMux I__4589 (
            .O(N__28308),
            .I(N__28260));
    LocalMux I__4588 (
            .O(N__28305),
            .I(N__28257));
    InMux I__4587 (
            .O(N__28304),
            .I(N__28254));
    InMux I__4586 (
            .O(N__28303),
            .I(N__28245));
    InMux I__4585 (
            .O(N__28302),
            .I(N__28245));
    InMux I__4584 (
            .O(N__28301),
            .I(N__28245));
    InMux I__4583 (
            .O(N__28300),
            .I(N__28245));
    LocalMux I__4582 (
            .O(N__28297),
            .I(N__28240));
    LocalMux I__4581 (
            .O(N__28290),
            .I(N__28240));
    InMux I__4580 (
            .O(N__28289),
            .I(N__28237));
    InMux I__4579 (
            .O(N__28288),
            .I(N__28230));
    InMux I__4578 (
            .O(N__28287),
            .I(N__28230));
    InMux I__4577 (
            .O(N__28286),
            .I(N__28230));
    InMux I__4576 (
            .O(N__28285),
            .I(N__28221));
    InMux I__4575 (
            .O(N__28284),
            .I(N__28221));
    InMux I__4574 (
            .O(N__28283),
            .I(N__28221));
    InMux I__4573 (
            .O(N__28282),
            .I(N__28221));
    InMux I__4572 (
            .O(N__28281),
            .I(N__28213));
    InMux I__4571 (
            .O(N__28278),
            .I(N__28213));
    InMux I__4570 (
            .O(N__28277),
            .I(N__28213));
    CascadeMux I__4569 (
            .O(N__28276),
            .I(N__28208));
    CascadeMux I__4568 (
            .O(N__28275),
            .I(N__28204));
    CascadeMux I__4567 (
            .O(N__28274),
            .I(N__28200));
    CascadeMux I__4566 (
            .O(N__28273),
            .I(N__28196));
    CascadeMux I__4565 (
            .O(N__28272),
            .I(N__28192));
    CascadeMux I__4564 (
            .O(N__28271),
            .I(N__28188));
    CascadeMux I__4563 (
            .O(N__28270),
            .I(N__28184));
    CascadeMux I__4562 (
            .O(N__28269),
            .I(N__28180));
    CascadeMux I__4561 (
            .O(N__28268),
            .I(N__28176));
    CascadeMux I__4560 (
            .O(N__28267),
            .I(N__28172));
    CascadeMux I__4559 (
            .O(N__28266),
            .I(N__28168));
    LocalMux I__4558 (
            .O(N__28263),
            .I(N__28161));
    LocalMux I__4557 (
            .O(N__28260),
            .I(N__28158));
    Span4Mux_s1_v I__4556 (
            .O(N__28257),
            .I(N__28153));
    LocalMux I__4555 (
            .O(N__28254),
            .I(N__28153));
    LocalMux I__4554 (
            .O(N__28245),
            .I(N__28150));
    Span4Mux_v I__4553 (
            .O(N__28240),
            .I(N__28141));
    LocalMux I__4552 (
            .O(N__28237),
            .I(N__28141));
    LocalMux I__4551 (
            .O(N__28230),
            .I(N__28141));
    LocalMux I__4550 (
            .O(N__28221),
            .I(N__28141));
    InMux I__4549 (
            .O(N__28220),
            .I(N__28138));
    LocalMux I__4548 (
            .O(N__28213),
            .I(N__28135));
    InMux I__4547 (
            .O(N__28212),
            .I(N__28132));
    InMux I__4546 (
            .O(N__28211),
            .I(N__28117));
    InMux I__4545 (
            .O(N__28208),
            .I(N__28117));
    InMux I__4544 (
            .O(N__28207),
            .I(N__28117));
    InMux I__4543 (
            .O(N__28204),
            .I(N__28117));
    InMux I__4542 (
            .O(N__28203),
            .I(N__28117));
    InMux I__4541 (
            .O(N__28200),
            .I(N__28117));
    InMux I__4540 (
            .O(N__28199),
            .I(N__28117));
    InMux I__4539 (
            .O(N__28196),
            .I(N__28100));
    InMux I__4538 (
            .O(N__28195),
            .I(N__28100));
    InMux I__4537 (
            .O(N__28192),
            .I(N__28100));
    InMux I__4536 (
            .O(N__28191),
            .I(N__28100));
    InMux I__4535 (
            .O(N__28188),
            .I(N__28100));
    InMux I__4534 (
            .O(N__28187),
            .I(N__28100));
    InMux I__4533 (
            .O(N__28184),
            .I(N__28100));
    InMux I__4532 (
            .O(N__28183),
            .I(N__28100));
    InMux I__4531 (
            .O(N__28180),
            .I(N__28083));
    InMux I__4530 (
            .O(N__28179),
            .I(N__28083));
    InMux I__4529 (
            .O(N__28176),
            .I(N__28083));
    InMux I__4528 (
            .O(N__28175),
            .I(N__28083));
    InMux I__4527 (
            .O(N__28172),
            .I(N__28083));
    InMux I__4526 (
            .O(N__28171),
            .I(N__28083));
    InMux I__4525 (
            .O(N__28168),
            .I(N__28083));
    InMux I__4524 (
            .O(N__28167),
            .I(N__28083));
    CascadeMux I__4523 (
            .O(N__28166),
            .I(N__28079));
    CascadeMux I__4522 (
            .O(N__28165),
            .I(N__28075));
    CascadeMux I__4521 (
            .O(N__28164),
            .I(N__28071));
    Span12Mux_v I__4520 (
            .O(N__28161),
            .I(N__28067));
    Span12Mux_s1_h I__4519 (
            .O(N__28158),
            .I(N__28062));
    Sp12to4 I__4518 (
            .O(N__28153),
            .I(N__28062));
    Sp12to4 I__4517 (
            .O(N__28150),
            .I(N__28057));
    Sp12to4 I__4516 (
            .O(N__28141),
            .I(N__28057));
    LocalMux I__4515 (
            .O(N__28138),
            .I(N__28054));
    Span4Mux_h I__4514 (
            .O(N__28135),
            .I(N__28051));
    LocalMux I__4513 (
            .O(N__28132),
            .I(N__28048));
    LocalMux I__4512 (
            .O(N__28117),
            .I(N__28041));
    LocalMux I__4511 (
            .O(N__28100),
            .I(N__28041));
    LocalMux I__4510 (
            .O(N__28083),
            .I(N__28041));
    InMux I__4509 (
            .O(N__28082),
            .I(N__28026));
    InMux I__4508 (
            .O(N__28079),
            .I(N__28026));
    InMux I__4507 (
            .O(N__28078),
            .I(N__28026));
    InMux I__4506 (
            .O(N__28075),
            .I(N__28026));
    InMux I__4505 (
            .O(N__28074),
            .I(N__28026));
    InMux I__4504 (
            .O(N__28071),
            .I(N__28026));
    InMux I__4503 (
            .O(N__28070),
            .I(N__28026));
    Span12Mux_h I__4502 (
            .O(N__28067),
            .I(N__28019));
    Span12Mux_v I__4501 (
            .O(N__28062),
            .I(N__28019));
    Span12Mux_v I__4500 (
            .O(N__28057),
            .I(N__28019));
    Span4Mux_v I__4499 (
            .O(N__28054),
            .I(N__28016));
    Span4Mux_v I__4498 (
            .O(N__28051),
            .I(N__28007));
    Span4Mux_v I__4497 (
            .O(N__28048),
            .I(N__28007));
    Span4Mux_v I__4496 (
            .O(N__28041),
            .I(N__28007));
    LocalMux I__4495 (
            .O(N__28026),
            .I(N__28007));
    Odrv12 I__4494 (
            .O(N__28019),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4493 (
            .O(N__28016),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4492 (
            .O(N__28007),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__4491 (
            .O(N__28000),
            .I(N__27997));
    InMux I__4490 (
            .O(N__27997),
            .I(N__27992));
    CascadeMux I__4489 (
            .O(N__27996),
            .I(N__27987));
    InMux I__4488 (
            .O(N__27995),
            .I(N__27984));
    LocalMux I__4487 (
            .O(N__27992),
            .I(N__27981));
    InMux I__4486 (
            .O(N__27991),
            .I(N__27976));
    InMux I__4485 (
            .O(N__27990),
            .I(N__27976));
    InMux I__4484 (
            .O(N__27987),
            .I(N__27973));
    LocalMux I__4483 (
            .O(N__27984),
            .I(N__27969));
    Span4Mux_h I__4482 (
            .O(N__27981),
            .I(N__27964));
    LocalMux I__4481 (
            .O(N__27976),
            .I(N__27964));
    LocalMux I__4480 (
            .O(N__27973),
            .I(N__27961));
    InMux I__4479 (
            .O(N__27972),
            .I(N__27958));
    Span4Mux_h I__4478 (
            .O(N__27969),
            .I(N__27955));
    Span4Mux_v I__4477 (
            .O(N__27964),
            .I(N__27952));
    Odrv4 I__4476 (
            .O(N__27961),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__4475 (
            .O(N__27958),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__4474 (
            .O(N__27955),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__4473 (
            .O(N__27952),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__4472 (
            .O(N__27943),
            .I(N__27939));
    CascadeMux I__4471 (
            .O(N__27942),
            .I(N__27936));
    LocalMux I__4470 (
            .O(N__27939),
            .I(N__27933));
    InMux I__4469 (
            .O(N__27936),
            .I(N__27930));
    Odrv12 I__4468 (
            .O(N__27933),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    LocalMux I__4467 (
            .O(N__27930),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    InMux I__4466 (
            .O(N__27925),
            .I(N__27921));
    InMux I__4465 (
            .O(N__27924),
            .I(N__27918));
    LocalMux I__4464 (
            .O(N__27921),
            .I(N__27915));
    LocalMux I__4463 (
            .O(N__27918),
            .I(N__27912));
    Span4Mux_v I__4462 (
            .O(N__27915),
            .I(N__27907));
    Span4Mux_h I__4461 (
            .O(N__27912),
            .I(N__27907));
    Odrv4 I__4460 (
            .O(N__27907),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    CascadeMux I__4459 (
            .O(N__27904),
            .I(N__27901));
    InMux I__4458 (
            .O(N__27901),
            .I(N__27898));
    LocalMux I__4457 (
            .O(N__27898),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__4456 (
            .O(N__27895),
            .I(N__27892));
    LocalMux I__4455 (
            .O(N__27892),
            .I(N__27888));
    InMux I__4454 (
            .O(N__27891),
            .I(N__27885));
    Span4Mux_h I__4453 (
            .O(N__27888),
            .I(N__27882));
    LocalMux I__4452 (
            .O(N__27885),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__4451 (
            .O(N__27882),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__4450 (
            .O(N__27877),
            .I(N__27874));
    LocalMux I__4449 (
            .O(N__27874),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    CascadeMux I__4448 (
            .O(N__27871),
            .I(N__27868));
    InMux I__4447 (
            .O(N__27868),
            .I(N__27865));
    LocalMux I__4446 (
            .O(N__27865),
            .I(N__27862));
    Span4Mux_v I__4445 (
            .O(N__27862),
            .I(N__27859));
    Odrv4 I__4444 (
            .O(N__27859),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__4443 (
            .O(N__27856),
            .I(N__27853));
    LocalMux I__4442 (
            .O(N__27853),
            .I(N__27850));
    Span4Mux_v I__4441 (
            .O(N__27850),
            .I(N__27847));
    Odrv4 I__4440 (
            .O(N__27847),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__4439 (
            .O(N__27844),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__4438 (
            .O(N__27841),
            .I(N__27838));
    LocalMux I__4437 (
            .O(N__27838),
            .I(N__27835));
    Span4Mux_v I__4436 (
            .O(N__27835),
            .I(N__27832));
    Odrv4 I__4435 (
            .O(N__27832),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__4434 (
            .O(N__27829),
            .I(N__27826));
    LocalMux I__4433 (
            .O(N__27826),
            .I(N__27823));
    Odrv12 I__4432 (
            .O(N__27823),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__4431 (
            .O(N__27820),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    InMux I__4430 (
            .O(N__27817),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__4429 (
            .O(N__27814),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__4428 (
            .O(N__27811),
            .I(bfn_11_18_0_));
    InMux I__4427 (
            .O(N__27808),
            .I(N__27805));
    LocalMux I__4426 (
            .O(N__27805),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__4425 (
            .O(N__27802),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    CascadeMux I__4424 (
            .O(N__27799),
            .I(N__27796));
    InMux I__4423 (
            .O(N__27796),
            .I(N__27793));
    LocalMux I__4422 (
            .O(N__27793),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__4421 (
            .O(N__27790),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__4420 (
            .O(N__27787),
            .I(N__27784));
    LocalMux I__4419 (
            .O(N__27784),
            .I(N__27781));
    Odrv12 I__4418 (
            .O(N__27781),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__4417 (
            .O(N__27778),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__4416 (
            .O(N__27775),
            .I(N__27772));
    LocalMux I__4415 (
            .O(N__27772),
            .I(N__27769));
    Odrv12 I__4414 (
            .O(N__27769),
            .I(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ));
    CascadeMux I__4413 (
            .O(N__27766),
            .I(N__27763));
    InMux I__4412 (
            .O(N__27763),
            .I(N__27760));
    LocalMux I__4411 (
            .O(N__27760),
            .I(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ));
    InMux I__4410 (
            .O(N__27757),
            .I(N__27754));
    LocalMux I__4409 (
            .O(N__27754),
            .I(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ));
    CascadeMux I__4408 (
            .O(N__27751),
            .I(N__27748));
    InMux I__4407 (
            .O(N__27748),
            .I(N__27745));
    LocalMux I__4406 (
            .O(N__27745),
            .I(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ));
    InMux I__4405 (
            .O(N__27742),
            .I(N__27739));
    LocalMux I__4404 (
            .O(N__27739),
            .I(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ));
    CascadeMux I__4403 (
            .O(N__27736),
            .I(N__27733));
    InMux I__4402 (
            .O(N__27733),
            .I(N__27730));
    LocalMux I__4401 (
            .O(N__27730),
            .I(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ));
    CascadeMux I__4400 (
            .O(N__27727),
            .I(N__27724));
    InMux I__4399 (
            .O(N__27724),
            .I(N__27721));
    LocalMux I__4398 (
            .O(N__27721),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    CascadeMux I__4397 (
            .O(N__27718),
            .I(N__27715));
    InMux I__4396 (
            .O(N__27715),
            .I(N__27712));
    LocalMux I__4395 (
            .O(N__27712),
            .I(N__27709));
    Odrv4 I__4394 (
            .O(N__27709),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    CascadeMux I__4393 (
            .O(N__27706),
            .I(N__27703));
    InMux I__4392 (
            .O(N__27703),
            .I(N__27700));
    LocalMux I__4391 (
            .O(N__27700),
            .I(N__27697));
    Span4Mux_h I__4390 (
            .O(N__27697),
            .I(N__27694));
    Odrv4 I__4389 (
            .O(N__27694),
            .I(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ));
    InMux I__4388 (
            .O(N__27691),
            .I(N__27688));
    LocalMux I__4387 (
            .O(N__27688),
            .I(N__27685));
    Span4Mux_v I__4386 (
            .O(N__27685),
            .I(N__27682));
    Odrv4 I__4385 (
            .O(N__27682),
            .I(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ));
    CascadeMux I__4384 (
            .O(N__27679),
            .I(N__27676));
    InMux I__4383 (
            .O(N__27676),
            .I(N__27673));
    LocalMux I__4382 (
            .O(N__27673),
            .I(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ));
    InMux I__4381 (
            .O(N__27670),
            .I(N__27667));
    LocalMux I__4380 (
            .O(N__27667),
            .I(N__27663));
    InMux I__4379 (
            .O(N__27666),
            .I(N__27660));
    Span4Mux_v I__4378 (
            .O(N__27663),
            .I(N__27654));
    LocalMux I__4377 (
            .O(N__27660),
            .I(N__27654));
    InMux I__4376 (
            .O(N__27659),
            .I(N__27651));
    Span4Mux_h I__4375 (
            .O(N__27654),
            .I(N__27648));
    LocalMux I__4374 (
            .O(N__27651),
            .I(N__27645));
    Span4Mux_v I__4373 (
            .O(N__27648),
            .I(N__27642));
    Span4Mux_h I__4372 (
            .O(N__27645),
            .I(N__27639));
    Odrv4 I__4371 (
            .O(N__27642),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__4370 (
            .O(N__27639),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CEMux I__4369 (
            .O(N__27634),
            .I(N__27607));
    CEMux I__4368 (
            .O(N__27633),
            .I(N__27607));
    CEMux I__4367 (
            .O(N__27632),
            .I(N__27607));
    CEMux I__4366 (
            .O(N__27631),
            .I(N__27607));
    CEMux I__4365 (
            .O(N__27630),
            .I(N__27607));
    CEMux I__4364 (
            .O(N__27629),
            .I(N__27607));
    CEMux I__4363 (
            .O(N__27628),
            .I(N__27607));
    CEMux I__4362 (
            .O(N__27627),
            .I(N__27607));
    CEMux I__4361 (
            .O(N__27626),
            .I(N__27607));
    GlobalMux I__4360 (
            .O(N__27607),
            .I(N__27604));
    gio2CtrlBuf I__4359 (
            .O(N__27604),
            .I(\current_shift_inst.timer_s1.N_166_i_g ));
    InMux I__4358 (
            .O(N__27601),
            .I(N__27594));
    InMux I__4357 (
            .O(N__27600),
            .I(N__27594));
    InMux I__4356 (
            .O(N__27599),
            .I(N__27591));
    LocalMux I__4355 (
            .O(N__27594),
            .I(N__27588));
    LocalMux I__4354 (
            .O(N__27591),
            .I(N__27585));
    Span4Mux_h I__4353 (
            .O(N__27588),
            .I(N__27582));
    Span4Mux_v I__4352 (
            .O(N__27585),
            .I(N__27579));
    Odrv4 I__4351 (
            .O(N__27582),
            .I(\current_shift_inst.un4_control_input1_3 ));
    Odrv4 I__4350 (
            .O(N__27579),
            .I(\current_shift_inst.un4_control_input1_3 ));
    CascadeMux I__4349 (
            .O(N__27574),
            .I(N__27571));
    InMux I__4348 (
            .O(N__27571),
            .I(N__27565));
    InMux I__4347 (
            .O(N__27570),
            .I(N__27565));
    LocalMux I__4346 (
            .O(N__27565),
            .I(N__27562));
    Span4Mux_v I__4345 (
            .O(N__27562),
            .I(N__27559));
    Span4Mux_h I__4344 (
            .O(N__27559),
            .I(N__27554));
    InMux I__4343 (
            .O(N__27558),
            .I(N__27551));
    InMux I__4342 (
            .O(N__27557),
            .I(N__27548));
    Odrv4 I__4341 (
            .O(N__27554),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__4340 (
            .O(N__27551),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__4339 (
            .O(N__27548),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    CascadeMux I__4338 (
            .O(N__27541),
            .I(N__27538));
    InMux I__4337 (
            .O(N__27538),
            .I(N__27535));
    LocalMux I__4336 (
            .O(N__27535),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__4335 (
            .O(N__27532),
            .I(N__27529));
    LocalMux I__4334 (
            .O(N__27529),
            .I(N__27524));
    InMux I__4333 (
            .O(N__27528),
            .I(N__27521));
    CascadeMux I__4332 (
            .O(N__27527),
            .I(N__27518));
    Span4Mux_h I__4331 (
            .O(N__27524),
            .I(N__27515));
    LocalMux I__4330 (
            .O(N__27521),
            .I(N__27512));
    InMux I__4329 (
            .O(N__27518),
            .I(N__27509));
    Odrv4 I__4328 (
            .O(N__27515),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv4 I__4327 (
            .O(N__27512),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__4326 (
            .O(N__27509),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__4325 (
            .O(N__27502),
            .I(N__27499));
    LocalMux I__4324 (
            .O(N__27499),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__4323 (
            .O(N__27496),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__4322 (
            .O(N__27493),
            .I(N__27487));
    InMux I__4321 (
            .O(N__27492),
            .I(N__27487));
    LocalMux I__4320 (
            .O(N__27487),
            .I(N__27482));
    InMux I__4319 (
            .O(N__27486),
            .I(N__27477));
    InMux I__4318 (
            .O(N__27485),
            .I(N__27477));
    Span4Mux_h I__4317 (
            .O(N__27482),
            .I(N__27474));
    LocalMux I__4316 (
            .O(N__27477),
            .I(N__27471));
    Span4Mux_v I__4315 (
            .O(N__27474),
            .I(N__27468));
    Span12Mux_v I__4314 (
            .O(N__27471),
            .I(N__27465));
    Odrv4 I__4313 (
            .O(N__27468),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    Odrv12 I__4312 (
            .O(N__27465),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__4311 (
            .O(N__27460),
            .I(N__27457));
    InMux I__4310 (
            .O(N__27457),
            .I(N__27454));
    LocalMux I__4309 (
            .O(N__27454),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__4308 (
            .O(N__27451),
            .I(N__27448));
    InMux I__4307 (
            .O(N__27448),
            .I(N__27445));
    LocalMux I__4306 (
            .O(N__27445),
            .I(N__27442));
    Span4Mux_h I__4305 (
            .O(N__27442),
            .I(N__27439));
    Odrv4 I__4304 (
            .O(N__27439),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ));
    CascadeMux I__4303 (
            .O(N__27436),
            .I(N__27433));
    InMux I__4302 (
            .O(N__27433),
            .I(N__27429));
    InMux I__4301 (
            .O(N__27432),
            .I(N__27426));
    LocalMux I__4300 (
            .O(N__27429),
            .I(N__27423));
    LocalMux I__4299 (
            .O(N__27426),
            .I(N__27419));
    Span4Mux_v I__4298 (
            .O(N__27423),
            .I(N__27415));
    InMux I__4297 (
            .O(N__27422),
            .I(N__27412));
    Span4Mux_v I__4296 (
            .O(N__27419),
            .I(N__27409));
    InMux I__4295 (
            .O(N__27418),
            .I(N__27406));
    Span4Mux_h I__4294 (
            .O(N__27415),
            .I(N__27401));
    LocalMux I__4293 (
            .O(N__27412),
            .I(N__27401));
    Odrv4 I__4292 (
            .O(N__27409),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__4291 (
            .O(N__27406),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__4290 (
            .O(N__27401),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    InMux I__4289 (
            .O(N__27394),
            .I(N__27391));
    LocalMux I__4288 (
            .O(N__27391),
            .I(N__27388));
    Odrv4 I__4287 (
            .O(N__27388),
            .I(\current_shift_inst.PI_CTRL.integrator_i_23 ));
    InMux I__4286 (
            .O(N__27385),
            .I(N__27382));
    LocalMux I__4285 (
            .O(N__27382),
            .I(N__27379));
    Odrv4 I__4284 (
            .O(N__27379),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    CascadeMux I__4283 (
            .O(N__27376),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    InMux I__4282 (
            .O(N__27373),
            .I(N__27370));
    LocalMux I__4281 (
            .O(N__27370),
            .I(N__27367));
    Odrv4 I__4280 (
            .O(N__27367),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__4279 (
            .O(N__27364),
            .I(N__27361));
    LocalMux I__4278 (
            .O(N__27361),
            .I(N__27358));
    Span4Mux_h I__4277 (
            .O(N__27358),
            .I(N__27355));
    Odrv4 I__4276 (
            .O(N__27355),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    CascadeMux I__4275 (
            .O(N__27352),
            .I(N__27349));
    InMux I__4274 (
            .O(N__27349),
            .I(N__27345));
    InMux I__4273 (
            .O(N__27348),
            .I(N__27342));
    LocalMux I__4272 (
            .O(N__27345),
            .I(N__27339));
    LocalMux I__4271 (
            .O(N__27342),
            .I(N__27336));
    Span4Mux_v I__4270 (
            .O(N__27339),
            .I(N__27331));
    Span4Mux_v I__4269 (
            .O(N__27336),
            .I(N__27328));
    InMux I__4268 (
            .O(N__27335),
            .I(N__27325));
    InMux I__4267 (
            .O(N__27334),
            .I(N__27322));
    Span4Mux_v I__4266 (
            .O(N__27331),
            .I(N__27319));
    Span4Mux_h I__4265 (
            .O(N__27328),
            .I(N__27314));
    LocalMux I__4264 (
            .O(N__27325),
            .I(N__27314));
    LocalMux I__4263 (
            .O(N__27322),
            .I(N__27311));
    Odrv4 I__4262 (
            .O(N__27319),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__4261 (
            .O(N__27314),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv12 I__4260 (
            .O(N__27311),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__4259 (
            .O(N__27304),
            .I(N__27300));
    InMux I__4258 (
            .O(N__27303),
            .I(N__27296));
    LocalMux I__4257 (
            .O(N__27300),
            .I(N__27293));
    InMux I__4256 (
            .O(N__27299),
            .I(N__27290));
    LocalMux I__4255 (
            .O(N__27296),
            .I(N__27287));
    Odrv4 I__4254 (
            .O(N__27293),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__4253 (
            .O(N__27290),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv12 I__4252 (
            .O(N__27287),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__4251 (
            .O(N__27280),
            .I(N__27276));
    InMux I__4250 (
            .O(N__27279),
            .I(N__27273));
    LocalMux I__4249 (
            .O(N__27276),
            .I(N__27268));
    LocalMux I__4248 (
            .O(N__27273),
            .I(N__27268));
    Span4Mux_v I__4247 (
            .O(N__27268),
            .I(N__27263));
    InMux I__4246 (
            .O(N__27267),
            .I(N__27260));
    InMux I__4245 (
            .O(N__27266),
            .I(N__27257));
    Span4Mux_h I__4244 (
            .O(N__27263),
            .I(N__27252));
    LocalMux I__4243 (
            .O(N__27260),
            .I(N__27252));
    LocalMux I__4242 (
            .O(N__27257),
            .I(N__27249));
    Span4Mux_v I__4241 (
            .O(N__27252),
            .I(N__27246));
    Span4Mux_v I__4240 (
            .O(N__27249),
            .I(N__27243));
    Odrv4 I__4239 (
            .O(N__27246),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv4 I__4238 (
            .O(N__27243),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    CascadeMux I__4237 (
            .O(N__27238),
            .I(N__27235));
    InMux I__4236 (
            .O(N__27235),
            .I(N__27229));
    InMux I__4235 (
            .O(N__27234),
            .I(N__27229));
    LocalMux I__4234 (
            .O(N__27229),
            .I(N__27226));
    Span4Mux_v I__4233 (
            .O(N__27226),
            .I(N__27222));
    InMux I__4232 (
            .O(N__27225),
            .I(N__27219));
    Odrv4 I__4231 (
            .O(N__27222),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__4230 (
            .O(N__27219),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__4229 (
            .O(N__27214),
            .I(N__27211));
    LocalMux I__4228 (
            .O(N__27211),
            .I(N__27208));
    Odrv4 I__4227 (
            .O(N__27208),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__4226 (
            .O(N__27205),
            .I(bfn_11_10_0_));
    CascadeMux I__4225 (
            .O(N__27202),
            .I(N__27199));
    InMux I__4224 (
            .O(N__27199),
            .I(N__27196));
    LocalMux I__4223 (
            .O(N__27196),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    CascadeMux I__4222 (
            .O(N__27193),
            .I(N__27190));
    InMux I__4221 (
            .O(N__27190),
            .I(N__27186));
    InMux I__4220 (
            .O(N__27189),
            .I(N__27182));
    LocalMux I__4219 (
            .O(N__27186),
            .I(N__27179));
    InMux I__4218 (
            .O(N__27185),
            .I(N__27176));
    LocalMux I__4217 (
            .O(N__27182),
            .I(N__27172));
    Span4Mux_v I__4216 (
            .O(N__27179),
            .I(N__27167));
    LocalMux I__4215 (
            .O(N__27176),
            .I(N__27167));
    InMux I__4214 (
            .O(N__27175),
            .I(N__27164));
    Odrv4 I__4213 (
            .O(N__27172),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__4212 (
            .O(N__27167),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__4211 (
            .O(N__27164),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__4210 (
            .O(N__27157),
            .I(N__27154));
    InMux I__4209 (
            .O(N__27154),
            .I(N__27151));
    LocalMux I__4208 (
            .O(N__27151),
            .I(\current_shift_inst.PI_CTRL.integrator_i_29 ));
    InMux I__4207 (
            .O(N__27148),
            .I(N__27144));
    InMux I__4206 (
            .O(N__27147),
            .I(N__27141));
    LocalMux I__4205 (
            .O(N__27144),
            .I(N__27137));
    LocalMux I__4204 (
            .O(N__27141),
            .I(N__27134));
    InMux I__4203 (
            .O(N__27140),
            .I(N__27130));
    Span4Mux_v I__4202 (
            .O(N__27137),
            .I(N__27125));
    Span4Mux_v I__4201 (
            .O(N__27134),
            .I(N__27125));
    InMux I__4200 (
            .O(N__27133),
            .I(N__27122));
    LocalMux I__4199 (
            .O(N__27130),
            .I(N__27119));
    Odrv4 I__4198 (
            .O(N__27125),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__4197 (
            .O(N__27122),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__4196 (
            .O(N__27119),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    CascadeMux I__4195 (
            .O(N__27112),
            .I(N__27109));
    InMux I__4194 (
            .O(N__27109),
            .I(N__27106));
    LocalMux I__4193 (
            .O(N__27106),
            .I(\current_shift_inst.PI_CTRL.integrator_i_28 ));
    InMux I__4192 (
            .O(N__27103),
            .I(N__27100));
    LocalMux I__4191 (
            .O(N__27100),
            .I(N__27097));
    Odrv12 I__4190 (
            .O(N__27097),
            .I(\current_shift_inst.PI_CTRL.integrator_i_11 ));
    InMux I__4189 (
            .O(N__27094),
            .I(N__27089));
    InMux I__4188 (
            .O(N__27093),
            .I(N__27084));
    InMux I__4187 (
            .O(N__27092),
            .I(N__27084));
    LocalMux I__4186 (
            .O(N__27089),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ));
    LocalMux I__4185 (
            .O(N__27084),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ));
    InMux I__4184 (
            .O(N__27079),
            .I(N__27076));
    LocalMux I__4183 (
            .O(N__27076),
            .I(\current_shift_inst.PI_CTRL.integrator_i_25 ));
    InMux I__4182 (
            .O(N__27073),
            .I(N__27070));
    LocalMux I__4181 (
            .O(N__27070),
            .I(N__27067));
    Odrv4 I__4180 (
            .O(N__27067),
            .I(\current_shift_inst.PI_CTRL.integrator_i_26 ));
    InMux I__4179 (
            .O(N__27064),
            .I(N__27061));
    LocalMux I__4178 (
            .O(N__27061),
            .I(N__27058));
    Span4Mux_h I__4177 (
            .O(N__27058),
            .I(N__27055));
    Span4Mux_v I__4176 (
            .O(N__27055),
            .I(N__27052));
    Odrv4 I__4175 (
            .O(N__27052),
            .I(il_min_comp1_D1));
    InMux I__4174 (
            .O(N__27049),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ));
    InMux I__4173 (
            .O(N__27046),
            .I(N__27043));
    LocalMux I__4172 (
            .O(N__27043),
            .I(N__27040));
    Odrv4 I__4171 (
            .O(N__27040),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__4170 (
            .O(N__27037),
            .I(bfn_11_9_0_));
    CascadeMux I__4169 (
            .O(N__27034),
            .I(N__27031));
    InMux I__4168 (
            .O(N__27031),
            .I(N__27028));
    LocalMux I__4167 (
            .O(N__27028),
            .I(N__27025));
    Odrv4 I__4166 (
            .O(N__27025),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__4165 (
            .O(N__27022),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ));
    InMux I__4164 (
            .O(N__27019),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ));
    InMux I__4163 (
            .O(N__27016),
            .I(N__27013));
    LocalMux I__4162 (
            .O(N__27013),
            .I(N__27010));
    Odrv4 I__4161 (
            .O(N__27010),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__4160 (
            .O(N__27007),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ));
    CascadeMux I__4159 (
            .O(N__27004),
            .I(N__27001));
    InMux I__4158 (
            .O(N__27001),
            .I(N__26998));
    LocalMux I__4157 (
            .O(N__26998),
            .I(N__26995));
    Span4Mux_v I__4156 (
            .O(N__26995),
            .I(N__26992));
    Odrv4 I__4155 (
            .O(N__26992),
            .I(\current_shift_inst.PI_CTRL.integrator_i_27 ));
    InMux I__4154 (
            .O(N__26989),
            .I(N__26986));
    LocalMux I__4153 (
            .O(N__26986),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__4152 (
            .O(N__26983),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ));
    InMux I__4151 (
            .O(N__26980),
            .I(N__26977));
    LocalMux I__4150 (
            .O(N__26977),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__4149 (
            .O(N__26974),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ));
    InMux I__4148 (
            .O(N__26971),
            .I(N__26968));
    LocalMux I__4147 (
            .O(N__26968),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__4146 (
            .O(N__26965),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ));
    CascadeMux I__4145 (
            .O(N__26962),
            .I(N__26959));
    InMux I__4144 (
            .O(N__26959),
            .I(N__26956));
    LocalMux I__4143 (
            .O(N__26956),
            .I(N__26953));
    Span4Mux_h I__4142 (
            .O(N__26953),
            .I(N__26950));
    Odrv4 I__4141 (
            .O(N__26950),
            .I(\current_shift_inst.PI_CTRL.integrator_i_30 ));
    CascadeMux I__4140 (
            .O(N__26947),
            .I(N__26944));
    InMux I__4139 (
            .O(N__26944),
            .I(N__26941));
    LocalMux I__4138 (
            .O(N__26941),
            .I(N__26938));
    Odrv4 I__4137 (
            .O(N__26938),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__4136 (
            .O(N__26935),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ));
    InMux I__4135 (
            .O(N__26932),
            .I(N__26929));
    LocalMux I__4134 (
            .O(N__26929),
            .I(\current_shift_inst.PI_CTRL.integrator_i_14 ));
    CascadeMux I__4133 (
            .O(N__26926),
            .I(N__26923));
    InMux I__4132 (
            .O(N__26923),
            .I(N__26920));
    LocalMux I__4131 (
            .O(N__26920),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__4130 (
            .O(N__26917),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ));
    InMux I__4129 (
            .O(N__26914),
            .I(N__26911));
    LocalMux I__4128 (
            .O(N__26911),
            .I(N__26908));
    Odrv4 I__4127 (
            .O(N__26908),
            .I(\current_shift_inst.PI_CTRL.integrator_i_15 ));
    CascadeMux I__4126 (
            .O(N__26905),
            .I(N__26902));
    InMux I__4125 (
            .O(N__26902),
            .I(N__26899));
    LocalMux I__4124 (
            .O(N__26899),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__4123 (
            .O(N__26896),
            .I(bfn_11_8_0_));
    InMux I__4122 (
            .O(N__26893),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ));
    InMux I__4121 (
            .O(N__26890),
            .I(N__26887));
    LocalMux I__4120 (
            .O(N__26887),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__4119 (
            .O(N__26884),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ));
    InMux I__4118 (
            .O(N__26881),
            .I(N__26878));
    LocalMux I__4117 (
            .O(N__26878),
            .I(N__26875));
    Span4Mux_h I__4116 (
            .O(N__26875),
            .I(N__26872));
    Odrv4 I__4115 (
            .O(N__26872),
            .I(\current_shift_inst.PI_CTRL.integrator_i_18 ));
    CascadeMux I__4114 (
            .O(N__26869),
            .I(N__26866));
    InMux I__4113 (
            .O(N__26866),
            .I(N__26863));
    LocalMux I__4112 (
            .O(N__26863),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__4111 (
            .O(N__26860),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ));
    CascadeMux I__4110 (
            .O(N__26857),
            .I(N__26854));
    InMux I__4109 (
            .O(N__26854),
            .I(N__26851));
    LocalMux I__4108 (
            .O(N__26851),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__4107 (
            .O(N__26848),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ));
    InMux I__4106 (
            .O(N__26845),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ));
    InMux I__4105 (
            .O(N__26842),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ));
    CascadeMux I__4104 (
            .O(N__26839),
            .I(N__26836));
    InMux I__4103 (
            .O(N__26836),
            .I(N__26833));
    LocalMux I__4102 (
            .O(N__26833),
            .I(N__26830));
    Odrv12 I__4101 (
            .O(N__26830),
            .I(\current_shift_inst.PI_CTRL.integrator_i_22 ));
    CascadeMux I__4100 (
            .O(N__26827),
            .I(N__26824));
    InMux I__4099 (
            .O(N__26824),
            .I(N__26821));
    LocalMux I__4098 (
            .O(N__26821),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__4097 (
            .O(N__26818),
            .I(N__26815));
    LocalMux I__4096 (
            .O(N__26815),
            .I(N__26812));
    Span4Mux_h I__4095 (
            .O(N__26812),
            .I(N__26809));
    Odrv4 I__4094 (
            .O(N__26809),
            .I(\current_shift_inst.PI_CTRL.integrator_i_6 ));
    InMux I__4093 (
            .O(N__26806),
            .I(N__26803));
    LocalMux I__4092 (
            .O(N__26803),
            .I(N__26800));
    Odrv4 I__4091 (
            .O(N__26800),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__4090 (
            .O(N__26797),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ));
    InMux I__4089 (
            .O(N__26794),
            .I(N__26791));
    LocalMux I__4088 (
            .O(N__26791),
            .I(N__26788));
    Span4Mux_h I__4087 (
            .O(N__26788),
            .I(N__26785));
    Odrv4 I__4086 (
            .O(N__26785),
            .I(\current_shift_inst.PI_CTRL.integrator_i_7 ));
    InMux I__4085 (
            .O(N__26782),
            .I(bfn_11_7_0_));
    InMux I__4084 (
            .O(N__26779),
            .I(N__26776));
    LocalMux I__4083 (
            .O(N__26776),
            .I(N__26773));
    Odrv4 I__4082 (
            .O(N__26773),
            .I(\current_shift_inst.PI_CTRL.integrator_i_8 ));
    InMux I__4081 (
            .O(N__26770),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ));
    InMux I__4080 (
            .O(N__26767),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ));
    InMux I__4079 (
            .O(N__26764),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ));
    InMux I__4078 (
            .O(N__26761),
            .I(N__26758));
    LocalMux I__4077 (
            .O(N__26758),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__4076 (
            .O(N__26755),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ));
    InMux I__4075 (
            .O(N__26752),
            .I(N__26749));
    LocalMux I__4074 (
            .O(N__26749),
            .I(N__26746));
    Odrv4 I__4073 (
            .O(N__26746),
            .I(\current_shift_inst.PI_CTRL.integrator_i_12 ));
    CascadeMux I__4072 (
            .O(N__26743),
            .I(N__26740));
    InMux I__4071 (
            .O(N__26740),
            .I(N__26737));
    LocalMux I__4070 (
            .O(N__26737),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__4069 (
            .O(N__26734),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ));
    InMux I__4068 (
            .O(N__26731),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ));
    InMux I__4067 (
            .O(N__26728),
            .I(N__26725));
    LocalMux I__4066 (
            .O(N__26725),
            .I(N__26722));
    Odrv12 I__4065 (
            .O(N__26722),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ));
    InMux I__4064 (
            .O(N__26719),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ));
    InMux I__4063 (
            .O(N__26716),
            .I(N__26713));
    LocalMux I__4062 (
            .O(N__26713),
            .I(N__26710));
    Odrv4 I__4061 (
            .O(N__26710),
            .I(\current_shift_inst.PI_CTRL.integrator_i_1 ));
    InMux I__4060 (
            .O(N__26707),
            .I(N__26704));
    LocalMux I__4059 (
            .O(N__26704),
            .I(N__26701));
    Odrv4 I__4058 (
            .O(N__26701),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ));
    InMux I__4057 (
            .O(N__26698),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ));
    InMux I__4056 (
            .O(N__26695),
            .I(N__26692));
    LocalMux I__4055 (
            .O(N__26692),
            .I(\current_shift_inst.PI_CTRL.integrator_i_2 ));
    InMux I__4054 (
            .O(N__26689),
            .I(N__26686));
    LocalMux I__4053 (
            .O(N__26686),
            .I(N__26683));
    Odrv12 I__4052 (
            .O(N__26683),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__4051 (
            .O(N__26680),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ));
    InMux I__4050 (
            .O(N__26677),
            .I(N__26674));
    LocalMux I__4049 (
            .O(N__26674),
            .I(N__26671));
    Odrv4 I__4048 (
            .O(N__26671),
            .I(\current_shift_inst.PI_CTRL.integrator_i_3 ));
    CascadeMux I__4047 (
            .O(N__26668),
            .I(N__26665));
    InMux I__4046 (
            .O(N__26665),
            .I(N__26662));
    LocalMux I__4045 (
            .O(N__26662),
            .I(N__26659));
    Odrv4 I__4044 (
            .O(N__26659),
            .I(\current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7 ));
    InMux I__4043 (
            .O(N__26656),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ));
    InMux I__4042 (
            .O(N__26653),
            .I(N__26650));
    LocalMux I__4041 (
            .O(N__26650),
            .I(\current_shift_inst.PI_CTRL.integrator_i_4 ));
    InMux I__4040 (
            .O(N__26647),
            .I(N__26644));
    LocalMux I__4039 (
            .O(N__26644),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__4038 (
            .O(N__26641),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ));
    CascadeMux I__4037 (
            .O(N__26638),
            .I(N__26635));
    InMux I__4036 (
            .O(N__26635),
            .I(N__26632));
    LocalMux I__4035 (
            .O(N__26632),
            .I(\current_shift_inst.PI_CTRL.integrator_i_5 ));
    CascadeMux I__4034 (
            .O(N__26629),
            .I(N__26626));
    InMux I__4033 (
            .O(N__26626),
            .I(N__26623));
    LocalMux I__4032 (
            .O(N__26623),
            .I(N__26620));
    Odrv4 I__4031 (
            .O(N__26620),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__4030 (
            .O(N__26617),
            .I(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ));
    InMux I__4029 (
            .O(N__26614),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__4028 (
            .O(N__26611),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__4027 (
            .O(N__26608),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__4026 (
            .O(N__26605),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__4025 (
            .O(N__26602),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__4024 (
            .O(N__26599),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__4023 (
            .O(N__26596),
            .I(bfn_10_24_0_));
    InMux I__4022 (
            .O(N__26593),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__4021 (
            .O(N__26590),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__4020 (
            .O(N__26587),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__4019 (
            .O(N__26584),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__4018 (
            .O(N__26581),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__4017 (
            .O(N__26578),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__4016 (
            .O(N__26575),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__4015 (
            .O(N__26572),
            .I(bfn_10_25_0_));
    InMux I__4014 (
            .O(N__26569),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__4013 (
            .O(N__26566),
            .I(bfn_10_23_0_));
    InMux I__4012 (
            .O(N__26563),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__4011 (
            .O(N__26560),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__4010 (
            .O(N__26557),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__4009 (
            .O(N__26554),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__4008 (
            .O(N__26551),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__4007 (
            .O(N__26548),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__4006 (
            .O(N__26545),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__4005 (
            .O(N__26542),
            .I(N__26538));
    CascadeMux I__4004 (
            .O(N__26541),
            .I(N__26535));
    LocalMux I__4003 (
            .O(N__26538),
            .I(N__26532));
    InMux I__4002 (
            .O(N__26535),
            .I(N__26529));
    Span4Mux_v I__4001 (
            .O(N__26532),
            .I(N__26526));
    LocalMux I__4000 (
            .O(N__26529),
            .I(N__26523));
    Span4Mux_v I__3999 (
            .O(N__26526),
            .I(N__26520));
    Span4Mux_v I__3998 (
            .O(N__26523),
            .I(N__26517));
    Odrv4 I__3997 (
            .O(N__26520),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv4 I__3996 (
            .O(N__26517),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__3995 (
            .O(N__26512),
            .I(N__26509));
    LocalMux I__3994 (
            .O(N__26509),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    InMux I__3993 (
            .O(N__26506),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__3992 (
            .O(N__26503),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__3991 (
            .O(N__26500),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__3990 (
            .O(N__26497),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__3989 (
            .O(N__26494),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__3988 (
            .O(N__26491),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    CascadeMux I__3987 (
            .O(N__26488),
            .I(N__26485));
    InMux I__3986 (
            .O(N__26485),
            .I(N__26482));
    LocalMux I__3985 (
            .O(N__26482),
            .I(N__26478));
    CascadeMux I__3984 (
            .O(N__26481),
            .I(N__26475));
    Span4Mux_h I__3983 (
            .O(N__26478),
            .I(N__26470));
    InMux I__3982 (
            .O(N__26475),
            .I(N__26467));
    InMux I__3981 (
            .O(N__26474),
            .I(N__26464));
    InMux I__3980 (
            .O(N__26473),
            .I(N__26461));
    Span4Mux_h I__3979 (
            .O(N__26470),
            .I(N__26456));
    LocalMux I__3978 (
            .O(N__26467),
            .I(N__26456));
    LocalMux I__3977 (
            .O(N__26464),
            .I(N__26451));
    LocalMux I__3976 (
            .O(N__26461),
            .I(N__26451));
    Odrv4 I__3975 (
            .O(N__26456),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    Odrv12 I__3974 (
            .O(N__26451),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__3973 (
            .O(N__26446),
            .I(N__26443));
    LocalMux I__3972 (
            .O(N__26443),
            .I(N__26439));
    InMux I__3971 (
            .O(N__26442),
            .I(N__26435));
    Span4Mux_h I__3970 (
            .O(N__26439),
            .I(N__26432));
    InMux I__3969 (
            .O(N__26438),
            .I(N__26429));
    LocalMux I__3968 (
            .O(N__26435),
            .I(N__26426));
    Odrv4 I__3967 (
            .O(N__26432),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__3966 (
            .O(N__26429),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__3965 (
            .O(N__26426),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__3964 (
            .O(N__26419),
            .I(N__26416));
    LocalMux I__3963 (
            .O(N__26416),
            .I(N__26412));
    InMux I__3962 (
            .O(N__26415),
            .I(N__26409));
    Span4Mux_h I__3961 (
            .O(N__26412),
            .I(N__26406));
    LocalMux I__3960 (
            .O(N__26409),
            .I(N__26403));
    Odrv4 I__3959 (
            .O(N__26406),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv4 I__3958 (
            .O(N__26403),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__3957 (
            .O(N__26398),
            .I(N__26395));
    InMux I__3956 (
            .O(N__26395),
            .I(N__26392));
    LocalMux I__3955 (
            .O(N__26392),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    CascadeMux I__3954 (
            .O(N__26389),
            .I(N__26386));
    InMux I__3953 (
            .O(N__26386),
            .I(N__26383));
    LocalMux I__3952 (
            .O(N__26383),
            .I(N__26380));
    Odrv4 I__3951 (
            .O(N__26380),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__3950 (
            .O(N__26377),
            .I(N__26373));
    InMux I__3949 (
            .O(N__26376),
            .I(N__26370));
    LocalMux I__3948 (
            .O(N__26373),
            .I(N__26365));
    LocalMux I__3947 (
            .O(N__26370),
            .I(N__26362));
    InMux I__3946 (
            .O(N__26369),
            .I(N__26359));
    InMux I__3945 (
            .O(N__26368),
            .I(N__26356));
    Span4Mux_h I__3944 (
            .O(N__26365),
            .I(N__26349));
    Span4Mux_v I__3943 (
            .O(N__26362),
            .I(N__26349));
    LocalMux I__3942 (
            .O(N__26359),
            .I(N__26349));
    LocalMux I__3941 (
            .O(N__26356),
            .I(N__26346));
    Odrv4 I__3940 (
            .O(N__26349),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv12 I__3939 (
            .O(N__26346),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__3938 (
            .O(N__26341),
            .I(N__26338));
    LocalMux I__3937 (
            .O(N__26338),
            .I(N__26334));
    InMux I__3936 (
            .O(N__26337),
            .I(N__26331));
    Span4Mux_h I__3935 (
            .O(N__26334),
            .I(N__26325));
    LocalMux I__3934 (
            .O(N__26331),
            .I(N__26325));
    InMux I__3933 (
            .O(N__26330),
            .I(N__26322));
    Span4Mux_v I__3932 (
            .O(N__26325),
            .I(N__26319));
    LocalMux I__3931 (
            .O(N__26322),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__3930 (
            .O(N__26319),
            .I(\current_shift_inst.un4_control_input1_26 ));
    CascadeMux I__3929 (
            .O(N__26314),
            .I(N__26311));
    InMux I__3928 (
            .O(N__26311),
            .I(N__26307));
    InMux I__3927 (
            .O(N__26310),
            .I(N__26304));
    LocalMux I__3926 (
            .O(N__26307),
            .I(N__26299));
    LocalMux I__3925 (
            .O(N__26304),
            .I(N__26296));
    InMux I__3924 (
            .O(N__26303),
            .I(N__26293));
    InMux I__3923 (
            .O(N__26302),
            .I(N__26290));
    Span4Mux_v I__3922 (
            .O(N__26299),
            .I(N__26287));
    Span4Mux_h I__3921 (
            .O(N__26296),
            .I(N__26282));
    LocalMux I__3920 (
            .O(N__26293),
            .I(N__26282));
    LocalMux I__3919 (
            .O(N__26290),
            .I(N__26279));
    Odrv4 I__3918 (
            .O(N__26287),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv4 I__3917 (
            .O(N__26282),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    Odrv12 I__3916 (
            .O(N__26279),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    CascadeMux I__3915 (
            .O(N__26272),
            .I(N__26269));
    InMux I__3914 (
            .O(N__26269),
            .I(N__26266));
    LocalMux I__3913 (
            .O(N__26266),
            .I(N__26262));
    InMux I__3912 (
            .O(N__26265),
            .I(N__26259));
    Span4Mux_v I__3911 (
            .O(N__26262),
            .I(N__26255));
    LocalMux I__3910 (
            .O(N__26259),
            .I(N__26252));
    InMux I__3909 (
            .O(N__26258),
            .I(N__26249));
    Span4Mux_h I__3908 (
            .O(N__26255),
            .I(N__26244));
    Span4Mux_v I__3907 (
            .O(N__26252),
            .I(N__26244));
    LocalMux I__3906 (
            .O(N__26249),
            .I(N__26241));
    Odrv4 I__3905 (
            .O(N__26244),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv12 I__3904 (
            .O(N__26241),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CascadeMux I__3903 (
            .O(N__26236),
            .I(N__26233));
    InMux I__3902 (
            .O(N__26233),
            .I(N__26230));
    LocalMux I__3901 (
            .O(N__26230),
            .I(N__26227));
    Odrv12 I__3900 (
            .O(N__26227),
            .I(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ));
    InMux I__3899 (
            .O(N__26224),
            .I(N__26220));
    InMux I__3898 (
            .O(N__26223),
            .I(N__26217));
    LocalMux I__3897 (
            .O(N__26220),
            .I(N__26214));
    LocalMux I__3896 (
            .O(N__26217),
            .I(N__26211));
    Span4Mux_v I__3895 (
            .O(N__26214),
            .I(N__26208));
    Span4Mux_v I__3894 (
            .O(N__26211),
            .I(N__26203));
    Span4Mux_h I__3893 (
            .O(N__26208),
            .I(N__26200));
    InMux I__3892 (
            .O(N__26207),
            .I(N__26195));
    InMux I__3891 (
            .O(N__26206),
            .I(N__26195));
    Span4Mux_h I__3890 (
            .O(N__26203),
            .I(N__26190));
    Span4Mux_v I__3889 (
            .O(N__26200),
            .I(N__26190));
    LocalMux I__3888 (
            .O(N__26195),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__3887 (
            .O(N__26190),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__3886 (
            .O(N__26185),
            .I(N__26182));
    LocalMux I__3885 (
            .O(N__26182),
            .I(N__26177));
    InMux I__3884 (
            .O(N__26181),
            .I(N__26174));
    InMux I__3883 (
            .O(N__26180),
            .I(N__26171));
    Sp12to4 I__3882 (
            .O(N__26177),
            .I(N__26164));
    LocalMux I__3881 (
            .O(N__26174),
            .I(N__26164));
    LocalMux I__3880 (
            .O(N__26171),
            .I(N__26164));
    Span12Mux_v I__3879 (
            .O(N__26164),
            .I(N__26161));
    Odrv12 I__3878 (
            .O(N__26161),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    IoInMux I__3877 (
            .O(N__26158),
            .I(N__26155));
    LocalMux I__3876 (
            .O(N__26155),
            .I(N__26152));
    Span4Mux_s3_v I__3875 (
            .O(N__26152),
            .I(N__26149));
    Span4Mux_h I__3874 (
            .O(N__26149),
            .I(N__26146));
    Span4Mux_v I__3873 (
            .O(N__26146),
            .I(N__26143));
    Odrv4 I__3872 (
            .O(N__26143),
            .I(\delay_measurement_inst.delay_hc_timer.N_397_i ));
    InMux I__3871 (
            .O(N__26140),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    CascadeMux I__3870 (
            .O(N__26137),
            .I(N__26134));
    InMux I__3869 (
            .O(N__26134),
            .I(N__26129));
    InMux I__3868 (
            .O(N__26133),
            .I(N__26126));
    InMux I__3867 (
            .O(N__26132),
            .I(N__26123));
    LocalMux I__3866 (
            .O(N__26129),
            .I(N__26118));
    LocalMux I__3865 (
            .O(N__26126),
            .I(N__26118));
    LocalMux I__3864 (
            .O(N__26123),
            .I(N__26113));
    Span4Mux_v I__3863 (
            .O(N__26118),
            .I(N__26113));
    Span4Mux_v I__3862 (
            .O(N__26113),
            .I(N__26109));
    InMux I__3861 (
            .O(N__26112),
            .I(N__26106));
    Odrv4 I__3860 (
            .O(N__26109),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__3859 (
            .O(N__26106),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__3858 (
            .O(N__26101),
            .I(N__26098));
    LocalMux I__3857 (
            .O(N__26098),
            .I(N__26095));
    Span4Mux_h I__3856 (
            .O(N__26095),
            .I(N__26090));
    InMux I__3855 (
            .O(N__26094),
            .I(N__26087));
    InMux I__3854 (
            .O(N__26093),
            .I(N__26084));
    Odrv4 I__3853 (
            .O(N__26090),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__3852 (
            .O(N__26087),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__3851 (
            .O(N__26084),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__3850 (
            .O(N__26077),
            .I(N__26073));
    InMux I__3849 (
            .O(N__26076),
            .I(N__26070));
    InMux I__3848 (
            .O(N__26073),
            .I(N__26067));
    LocalMux I__3847 (
            .O(N__26070),
            .I(N__26060));
    LocalMux I__3846 (
            .O(N__26067),
            .I(N__26060));
    InMux I__3845 (
            .O(N__26066),
            .I(N__26057));
    InMux I__3844 (
            .O(N__26065),
            .I(N__26054));
    Span4Mux_v I__3843 (
            .O(N__26060),
            .I(N__26051));
    LocalMux I__3842 (
            .O(N__26057),
            .I(N__26048));
    LocalMux I__3841 (
            .O(N__26054),
            .I(N__26045));
    Span4Mux_v I__3840 (
            .O(N__26051),
            .I(N__26042));
    Span4Mux_h I__3839 (
            .O(N__26048),
            .I(N__26037));
    Span4Mux_v I__3838 (
            .O(N__26045),
            .I(N__26037));
    Odrv4 I__3837 (
            .O(N__26042),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__3836 (
            .O(N__26037),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__3835 (
            .O(N__26032),
            .I(N__26029));
    LocalMux I__3834 (
            .O(N__26029),
            .I(N__26025));
    InMux I__3833 (
            .O(N__26028),
            .I(N__26022));
    Span4Mux_v I__3832 (
            .O(N__26025),
            .I(N__26018));
    LocalMux I__3831 (
            .O(N__26022),
            .I(N__26015));
    InMux I__3830 (
            .O(N__26021),
            .I(N__26012));
    Span4Mux_h I__3829 (
            .O(N__26018),
            .I(N__26009));
    Span4Mux_v I__3828 (
            .O(N__26015),
            .I(N__26006));
    LocalMux I__3827 (
            .O(N__26012),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__3826 (
            .O(N__26009),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__3825 (
            .O(N__26006),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__3824 (
            .O(N__25999),
            .I(N__25996));
    LocalMux I__3823 (
            .O(N__25996),
            .I(N__25991));
    InMux I__3822 (
            .O(N__25995),
            .I(N__25988));
    InMux I__3821 (
            .O(N__25994),
            .I(N__25985));
    Span4Mux_h I__3820 (
            .O(N__25991),
            .I(N__25980));
    LocalMux I__3819 (
            .O(N__25988),
            .I(N__25980));
    LocalMux I__3818 (
            .O(N__25985),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__3817 (
            .O(N__25980),
            .I(\current_shift_inst.un4_control_input1_16 ));
    CascadeMux I__3816 (
            .O(N__25975),
            .I(N__25972));
    InMux I__3815 (
            .O(N__25972),
            .I(N__25968));
    CascadeMux I__3814 (
            .O(N__25971),
            .I(N__25965));
    LocalMux I__3813 (
            .O(N__25968),
            .I(N__25962));
    InMux I__3812 (
            .O(N__25965),
            .I(N__25959));
    Span4Mux_v I__3811 (
            .O(N__25962),
            .I(N__25953));
    LocalMux I__3810 (
            .O(N__25959),
            .I(N__25953));
    InMux I__3809 (
            .O(N__25958),
            .I(N__25949));
    Span4Mux_h I__3808 (
            .O(N__25953),
            .I(N__25946));
    InMux I__3807 (
            .O(N__25952),
            .I(N__25943));
    LocalMux I__3806 (
            .O(N__25949),
            .I(N__25940));
    Span4Mux_v I__3805 (
            .O(N__25946),
            .I(N__25937));
    LocalMux I__3804 (
            .O(N__25943),
            .I(N__25934));
    Span4Mux_v I__3803 (
            .O(N__25940),
            .I(N__25931));
    Odrv4 I__3802 (
            .O(N__25937),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__3801 (
            .O(N__25934),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__3800 (
            .O(N__25931),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__3799 (
            .O(N__25924),
            .I(N__25919));
    InMux I__3798 (
            .O(N__25923),
            .I(N__25916));
    InMux I__3797 (
            .O(N__25922),
            .I(N__25912));
    LocalMux I__3796 (
            .O(N__25919),
            .I(N__25909));
    LocalMux I__3795 (
            .O(N__25916),
            .I(N__25906));
    InMux I__3794 (
            .O(N__25915),
            .I(N__25903));
    LocalMux I__3793 (
            .O(N__25912),
            .I(N__25900));
    Span4Mux_h I__3792 (
            .O(N__25909),
            .I(N__25897));
    Span12Mux_v I__3791 (
            .O(N__25906),
            .I(N__25894));
    LocalMux I__3790 (
            .O(N__25903),
            .I(N__25891));
    Span4Mux_v I__3789 (
            .O(N__25900),
            .I(N__25888));
    Odrv4 I__3788 (
            .O(N__25897),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv12 I__3787 (
            .O(N__25894),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__3786 (
            .O(N__25891),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__3785 (
            .O(N__25888),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    CascadeMux I__3784 (
            .O(N__25879),
            .I(N__25876));
    InMux I__3783 (
            .O(N__25876),
            .I(N__25872));
    InMux I__3782 (
            .O(N__25875),
            .I(N__25868));
    LocalMux I__3781 (
            .O(N__25872),
            .I(N__25865));
    InMux I__3780 (
            .O(N__25871),
            .I(N__25862));
    LocalMux I__3779 (
            .O(N__25868),
            .I(N__25859));
    Span4Mux_h I__3778 (
            .O(N__25865),
            .I(N__25854));
    LocalMux I__3777 (
            .O(N__25862),
            .I(N__25854));
    Span4Mux_v I__3776 (
            .O(N__25859),
            .I(N__25851));
    Span4Mux_v I__3775 (
            .O(N__25854),
            .I(N__25848));
    Odrv4 I__3774 (
            .O(N__25851),
            .I(\current_shift_inst.un4_control_input1_9 ));
    Odrv4 I__3773 (
            .O(N__25848),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__3772 (
            .O(N__25843),
            .I(N__25840));
    LocalMux I__3771 (
            .O(N__25840),
            .I(N__25837));
    Span4Mux_h I__3770 (
            .O(N__25837),
            .I(N__25834));
    Odrv4 I__3769 (
            .O(N__25834),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__3768 (
            .O(N__25831),
            .I(N__25828));
    LocalMux I__3767 (
            .O(N__25828),
            .I(N__25822));
    InMux I__3766 (
            .O(N__25827),
            .I(N__25819));
    InMux I__3765 (
            .O(N__25826),
            .I(N__25816));
    InMux I__3764 (
            .O(N__25825),
            .I(N__25813));
    Span4Mux_h I__3763 (
            .O(N__25822),
            .I(N__25808));
    LocalMux I__3762 (
            .O(N__25819),
            .I(N__25808));
    LocalMux I__3761 (
            .O(N__25816),
            .I(N__25803));
    LocalMux I__3760 (
            .O(N__25813),
            .I(N__25803));
    Odrv4 I__3759 (
            .O(N__25808),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv12 I__3758 (
            .O(N__25803),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__3757 (
            .O(N__25798),
            .I(N__25795));
    LocalMux I__3756 (
            .O(N__25795),
            .I(N__25791));
    InMux I__3755 (
            .O(N__25794),
            .I(N__25787));
    Span4Mux_h I__3754 (
            .O(N__25791),
            .I(N__25784));
    InMux I__3753 (
            .O(N__25790),
            .I(N__25781));
    LocalMux I__3752 (
            .O(N__25787),
            .I(N__25778));
    Odrv4 I__3751 (
            .O(N__25784),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__3750 (
            .O(N__25781),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv12 I__3749 (
            .O(N__25778),
            .I(\current_shift_inst.un4_control_input1_27 ));
    CascadeMux I__3748 (
            .O(N__25771),
            .I(N__25768));
    InMux I__3747 (
            .O(N__25768),
            .I(N__25765));
    LocalMux I__3746 (
            .O(N__25765),
            .I(N__25762));
    Odrv4 I__3745 (
            .O(N__25762),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__3744 (
            .O(N__25759),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__3743 (
            .O(N__25756),
            .I(N__25753));
    LocalMux I__3742 (
            .O(N__25753),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__3741 (
            .O(N__25750),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    CascadeMux I__3740 (
            .O(N__25747),
            .I(N__25744));
    InMux I__3739 (
            .O(N__25744),
            .I(N__25741));
    LocalMux I__3738 (
            .O(N__25741),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__3737 (
            .O(N__25738),
            .I(bfn_10_16_0_));
    InMux I__3736 (
            .O(N__25735),
            .I(N__25732));
    LocalMux I__3735 (
            .O(N__25732),
            .I(N__25729));
    Odrv12 I__3734 (
            .O(N__25729),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__3733 (
            .O(N__25726),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    CascadeMux I__3732 (
            .O(N__25723),
            .I(N__25720));
    InMux I__3731 (
            .O(N__25720),
            .I(N__25717));
    LocalMux I__3730 (
            .O(N__25717),
            .I(N__25714));
    Odrv12 I__3729 (
            .O(N__25714),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__3728 (
            .O(N__25711),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__3727 (
            .O(N__25708),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    CascadeMux I__3726 (
            .O(N__25705),
            .I(N__25702));
    InMux I__3725 (
            .O(N__25702),
            .I(N__25699));
    LocalMux I__3724 (
            .O(N__25699),
            .I(N__25696));
    Odrv4 I__3723 (
            .O(N__25696),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__3722 (
            .O(N__25693),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__3721 (
            .O(N__25690),
            .I(N__25687));
    LocalMux I__3720 (
            .O(N__25687),
            .I(N__25684));
    Odrv4 I__3719 (
            .O(N__25684),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__3718 (
            .O(N__25681),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    CascadeMux I__3717 (
            .O(N__25678),
            .I(N__25675));
    InMux I__3716 (
            .O(N__25675),
            .I(N__25672));
    LocalMux I__3715 (
            .O(N__25672),
            .I(N__25669));
    Span4Mux_h I__3714 (
            .O(N__25669),
            .I(N__25666));
    Odrv4 I__3713 (
            .O(N__25666),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    InMux I__3712 (
            .O(N__25663),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    CascadeMux I__3711 (
            .O(N__25660),
            .I(N__25657));
    InMux I__3710 (
            .O(N__25657),
            .I(N__25654));
    LocalMux I__3709 (
            .O(N__25654),
            .I(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ));
    InMux I__3708 (
            .O(N__25651),
            .I(N__25648));
    LocalMux I__3707 (
            .O(N__25648),
            .I(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ));
    CascadeMux I__3706 (
            .O(N__25645),
            .I(N__25642));
    InMux I__3705 (
            .O(N__25642),
            .I(N__25639));
    LocalMux I__3704 (
            .O(N__25639),
            .I(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ));
    InMux I__3703 (
            .O(N__25636),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__3702 (
            .O(N__25633),
            .I(N__25630));
    LocalMux I__3701 (
            .O(N__25630),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__3700 (
            .O(N__25627),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__3699 (
            .O(N__25624),
            .I(N__25621));
    LocalMux I__3698 (
            .O(N__25621),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    CascadeMux I__3697 (
            .O(N__25618),
            .I(N__25615));
    InMux I__3696 (
            .O(N__25615),
            .I(N__25612));
    LocalMux I__3695 (
            .O(N__25612),
            .I(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ));
    InMux I__3694 (
            .O(N__25609),
            .I(N__25606));
    LocalMux I__3693 (
            .O(N__25606),
            .I(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ));
    CascadeMux I__3692 (
            .O(N__25603),
            .I(N__25600));
    InMux I__3691 (
            .O(N__25600),
            .I(N__25597));
    LocalMux I__3690 (
            .O(N__25597),
            .I(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ));
    InMux I__3689 (
            .O(N__25594),
            .I(N__25591));
    LocalMux I__3688 (
            .O(N__25591),
            .I(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ));
    CascadeMux I__3687 (
            .O(N__25588),
            .I(N__25585));
    InMux I__3686 (
            .O(N__25585),
            .I(N__25582));
    LocalMux I__3685 (
            .O(N__25582),
            .I(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ));
    InMux I__3684 (
            .O(N__25579),
            .I(N__25576));
    LocalMux I__3683 (
            .O(N__25576),
            .I(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ));
    CascadeMux I__3682 (
            .O(N__25573),
            .I(N__25570));
    InMux I__3681 (
            .O(N__25570),
            .I(N__25567));
    LocalMux I__3680 (
            .O(N__25567),
            .I(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ));
    InMux I__3679 (
            .O(N__25564),
            .I(N__25561));
    LocalMux I__3678 (
            .O(N__25561),
            .I(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ));
    CascadeMux I__3677 (
            .O(N__25558),
            .I(N__25547));
    CascadeMux I__3676 (
            .O(N__25557),
            .I(N__25543));
    CascadeMux I__3675 (
            .O(N__25556),
            .I(N__25539));
    CascadeMux I__3674 (
            .O(N__25555),
            .I(N__25535));
    CascadeMux I__3673 (
            .O(N__25554),
            .I(N__25532));
    CascadeMux I__3672 (
            .O(N__25553),
            .I(N__25528));
    CascadeMux I__3671 (
            .O(N__25552),
            .I(N__25524));
    CascadeMux I__3670 (
            .O(N__25551),
            .I(N__25520));
    InMux I__3669 (
            .O(N__25550),
            .I(N__25501));
    InMux I__3668 (
            .O(N__25547),
            .I(N__25501));
    InMux I__3667 (
            .O(N__25546),
            .I(N__25501));
    InMux I__3666 (
            .O(N__25543),
            .I(N__25501));
    InMux I__3665 (
            .O(N__25542),
            .I(N__25501));
    InMux I__3664 (
            .O(N__25539),
            .I(N__25501));
    InMux I__3663 (
            .O(N__25538),
            .I(N__25501));
    InMux I__3662 (
            .O(N__25535),
            .I(N__25501));
    InMux I__3661 (
            .O(N__25532),
            .I(N__25484));
    InMux I__3660 (
            .O(N__25531),
            .I(N__25484));
    InMux I__3659 (
            .O(N__25528),
            .I(N__25484));
    InMux I__3658 (
            .O(N__25527),
            .I(N__25484));
    InMux I__3657 (
            .O(N__25524),
            .I(N__25484));
    InMux I__3656 (
            .O(N__25523),
            .I(N__25484));
    InMux I__3655 (
            .O(N__25520),
            .I(N__25484));
    InMux I__3654 (
            .O(N__25519),
            .I(N__25484));
    CascadeMux I__3653 (
            .O(N__25518),
            .I(N__25481));
    LocalMux I__3652 (
            .O(N__25501),
            .I(N__25475));
    LocalMux I__3651 (
            .O(N__25484),
            .I(N__25475));
    InMux I__3650 (
            .O(N__25481),
            .I(N__25470));
    InMux I__3649 (
            .O(N__25480),
            .I(N__25470));
    Span4Mux_v I__3648 (
            .O(N__25475),
            .I(N__25467));
    LocalMux I__3647 (
            .O(N__25470),
            .I(N__25464));
    Odrv4 I__3646 (
            .O(N__25467),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    Odrv12 I__3645 (
            .O(N__25464),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__3644 (
            .O(N__25459),
            .I(N__25456));
    LocalMux I__3643 (
            .O(N__25456),
            .I(N__25453));
    Span4Mux_h I__3642 (
            .O(N__25453),
            .I(N__25450));
    Odrv4 I__3641 (
            .O(N__25450),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__3640 (
            .O(N__25447),
            .I(N__25444));
    InMux I__3639 (
            .O(N__25444),
            .I(N__25441));
    LocalMux I__3638 (
            .O(N__25441),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__3637 (
            .O(N__25438),
            .I(N__25435));
    LocalMux I__3636 (
            .O(N__25435),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    CascadeMux I__3635 (
            .O(N__25432),
            .I(N__25429));
    InMux I__3634 (
            .O(N__25429),
            .I(N__25426));
    LocalMux I__3633 (
            .O(N__25426),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    CascadeMux I__3632 (
            .O(N__25423),
            .I(N__25420));
    InMux I__3631 (
            .O(N__25420),
            .I(N__25417));
    LocalMux I__3630 (
            .O(N__25417),
            .I(N__25414));
    Odrv12 I__3629 (
            .O(N__25414),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__3628 (
            .O(N__25411),
            .I(N__25408));
    LocalMux I__3627 (
            .O(N__25408),
            .I(N__25405));
    Odrv4 I__3626 (
            .O(N__25405),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__3625 (
            .O(N__25402),
            .I(N__25399));
    LocalMux I__3624 (
            .O(N__25399),
            .I(N__25396));
    Odrv12 I__3623 (
            .O(N__25396),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__3622 (
            .O(N__25393),
            .I(N__25390));
    LocalMux I__3621 (
            .O(N__25390),
            .I(N__25387));
    Odrv12 I__3620 (
            .O(N__25387),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__3619 (
            .O(N__25384),
            .I(N__25381));
    LocalMux I__3618 (
            .O(N__25381),
            .I(N__25376));
    InMux I__3617 (
            .O(N__25380),
            .I(N__25372));
    CascadeMux I__3616 (
            .O(N__25379),
            .I(N__25369));
    Span4Mux_h I__3615 (
            .O(N__25376),
            .I(N__25366));
    InMux I__3614 (
            .O(N__25375),
            .I(N__25363));
    LocalMux I__3613 (
            .O(N__25372),
            .I(N__25360));
    InMux I__3612 (
            .O(N__25369),
            .I(N__25357));
    Span4Mux_v I__3611 (
            .O(N__25366),
            .I(N__25350));
    LocalMux I__3610 (
            .O(N__25363),
            .I(N__25350));
    Span4Mux_v I__3609 (
            .O(N__25360),
            .I(N__25350));
    LocalMux I__3608 (
            .O(N__25357),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__3607 (
            .O(N__25350),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__3606 (
            .O(N__25345),
            .I(N__25333));
    InMux I__3605 (
            .O(N__25344),
            .I(N__25333));
    InMux I__3604 (
            .O(N__25343),
            .I(N__25333));
    InMux I__3603 (
            .O(N__25342),
            .I(N__25333));
    LocalMux I__3602 (
            .O(N__25333),
            .I(N__25304));
    InMux I__3601 (
            .O(N__25332),
            .I(N__25295));
    InMux I__3600 (
            .O(N__25331),
            .I(N__25295));
    InMux I__3599 (
            .O(N__25330),
            .I(N__25295));
    InMux I__3598 (
            .O(N__25329),
            .I(N__25295));
    InMux I__3597 (
            .O(N__25328),
            .I(N__25286));
    InMux I__3596 (
            .O(N__25327),
            .I(N__25286));
    InMux I__3595 (
            .O(N__25326),
            .I(N__25286));
    InMux I__3594 (
            .O(N__25325),
            .I(N__25286));
    InMux I__3593 (
            .O(N__25324),
            .I(N__25277));
    InMux I__3592 (
            .O(N__25323),
            .I(N__25277));
    InMux I__3591 (
            .O(N__25322),
            .I(N__25277));
    InMux I__3590 (
            .O(N__25321),
            .I(N__25277));
    InMux I__3589 (
            .O(N__25320),
            .I(N__25272));
    InMux I__3588 (
            .O(N__25319),
            .I(N__25272));
    InMux I__3587 (
            .O(N__25318),
            .I(N__25263));
    InMux I__3586 (
            .O(N__25317),
            .I(N__25263));
    InMux I__3585 (
            .O(N__25316),
            .I(N__25263));
    InMux I__3584 (
            .O(N__25315),
            .I(N__25263));
    InMux I__3583 (
            .O(N__25314),
            .I(N__25254));
    InMux I__3582 (
            .O(N__25313),
            .I(N__25254));
    InMux I__3581 (
            .O(N__25312),
            .I(N__25254));
    InMux I__3580 (
            .O(N__25311),
            .I(N__25254));
    InMux I__3579 (
            .O(N__25310),
            .I(N__25245));
    InMux I__3578 (
            .O(N__25309),
            .I(N__25245));
    InMux I__3577 (
            .O(N__25308),
            .I(N__25245));
    InMux I__3576 (
            .O(N__25307),
            .I(N__25245));
    Span4Mux_h I__3575 (
            .O(N__25304),
            .I(N__25240));
    LocalMux I__3574 (
            .O(N__25295),
            .I(N__25240));
    LocalMux I__3573 (
            .O(N__25286),
            .I(N__25235));
    LocalMux I__3572 (
            .O(N__25277),
            .I(N__25235));
    LocalMux I__3571 (
            .O(N__25272),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__3570 (
            .O(N__25263),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__3569 (
            .O(N__25254),
            .I(\current_shift_inst.timer_s1.running_i ));
    LocalMux I__3568 (
            .O(N__25245),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__3567 (
            .O(N__25240),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__3566 (
            .O(N__25235),
            .I(\current_shift_inst.timer_s1.running_i ));
    IoInMux I__3565 (
            .O(N__25222),
            .I(N__25219));
    LocalMux I__3564 (
            .O(N__25219),
            .I(N__25216));
    Span4Mux_s2_v I__3563 (
            .O(N__25216),
            .I(N__25213));
    Odrv4 I__3562 (
            .O(N__25213),
            .I(s4_phy_c));
    InMux I__3561 (
            .O(N__25210),
            .I(N__25207));
    LocalMux I__3560 (
            .O(N__25207),
            .I(il_max_comp1_D1));
    CascadeMux I__3559 (
            .O(N__25204),
            .I(N__25201));
    InMux I__3558 (
            .O(N__25201),
            .I(N__25198));
    LocalMux I__3557 (
            .O(N__25198),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__3556 (
            .O(N__25195),
            .I(N__25192));
    LocalMux I__3555 (
            .O(N__25192),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__3554 (
            .O(N__25189),
            .I(N__25186));
    InMux I__3553 (
            .O(N__25186),
            .I(N__25183));
    LocalMux I__3552 (
            .O(N__25183),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__3551 (
            .O(N__25180),
            .I(N__25177));
    LocalMux I__3550 (
            .O(N__25177),
            .I(N__25174));
    Odrv4 I__3549 (
            .O(N__25174),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    CascadeMux I__3548 (
            .O(N__25171),
            .I(N__25168));
    InMux I__3547 (
            .O(N__25168),
            .I(N__25165));
    LocalMux I__3546 (
            .O(N__25165),
            .I(N__25162));
    Span4Mux_v I__3545 (
            .O(N__25162),
            .I(N__25159));
    Odrv4 I__3544 (
            .O(N__25159),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__3543 (
            .O(N__25156),
            .I(N__25153));
    LocalMux I__3542 (
            .O(N__25153),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__3541 (
            .O(N__25150),
            .I(N__25147));
    InMux I__3540 (
            .O(N__25147),
            .I(N__25144));
    LocalMux I__3539 (
            .O(N__25144),
            .I(N__25141));
    Span4Mux_v I__3538 (
            .O(N__25141),
            .I(N__25138));
    Odrv4 I__3537 (
            .O(N__25138),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__3536 (
            .O(N__25135),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    IoInMux I__3535 (
            .O(N__25132),
            .I(N__25129));
    LocalMux I__3534 (
            .O(N__25129),
            .I(N__25126));
    Span12Mux_s3_v I__3533 (
            .O(N__25126),
            .I(N__25123));
    Odrv12 I__3532 (
            .O(N__25123),
            .I(s3_phy_c));
    CascadeMux I__3531 (
            .O(N__25120),
            .I(N__25117));
    InMux I__3530 (
            .O(N__25117),
            .I(N__25114));
    LocalMux I__3529 (
            .O(N__25114),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    InMux I__3528 (
            .O(N__25111),
            .I(N__25108));
    LocalMux I__3527 (
            .O(N__25108),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__3526 (
            .O(N__25105),
            .I(N__25102));
    InMux I__3525 (
            .O(N__25102),
            .I(N__25099));
    LocalMux I__3524 (
            .O(N__25099),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__3523 (
            .O(N__25096),
            .I(N__25093));
    LocalMux I__3522 (
            .O(N__25093),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__3521 (
            .O(N__25090),
            .I(N__25087));
    LocalMux I__3520 (
            .O(N__25087),
            .I(N__25084));
    Odrv4 I__3519 (
            .O(N__25084),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__3518 (
            .O(N__25081),
            .I(N__25078));
    InMux I__3517 (
            .O(N__25078),
            .I(N__25075));
    LocalMux I__3516 (
            .O(N__25075),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__3515 (
            .O(N__25072),
            .I(N__25069));
    LocalMux I__3514 (
            .O(N__25069),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    CascadeMux I__3513 (
            .O(N__25066),
            .I(N__25063));
    InMux I__3512 (
            .O(N__25063),
            .I(N__25060));
    LocalMux I__3511 (
            .O(N__25060),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__3510 (
            .O(N__25057),
            .I(N__25054));
    LocalMux I__3509 (
            .O(N__25054),
            .I(N__25051));
    Odrv4 I__3508 (
            .O(N__25051),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__3507 (
            .O(N__25048),
            .I(N__25045));
    InMux I__3506 (
            .O(N__25045),
            .I(N__25042));
    LocalMux I__3505 (
            .O(N__25042),
            .I(N__25039));
    Odrv4 I__3504 (
            .O(N__25039),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    CascadeMux I__3503 (
            .O(N__25036),
            .I(N__25033));
    InMux I__3502 (
            .O(N__25033),
            .I(N__25030));
    LocalMux I__3501 (
            .O(N__25030),
            .I(N__25027));
    Odrv12 I__3500 (
            .O(N__25027),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__3499 (
            .O(N__25024),
            .I(N__25021));
    LocalMux I__3498 (
            .O(N__25021),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    InMux I__3497 (
            .O(N__25018),
            .I(N__25015));
    LocalMux I__3496 (
            .O(N__25015),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__3495 (
            .O(N__25012),
            .I(N__25009));
    InMux I__3494 (
            .O(N__25009),
            .I(N__25006));
    LocalMux I__3493 (
            .O(N__25006),
            .I(N__25003));
    Odrv4 I__3492 (
            .O(N__25003),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__3491 (
            .O(N__25000),
            .I(N__24997));
    LocalMux I__3490 (
            .O(N__24997),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    CascadeMux I__3489 (
            .O(N__24994),
            .I(N__24991));
    InMux I__3488 (
            .O(N__24991),
            .I(N__24988));
    LocalMux I__3487 (
            .O(N__24988),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__3486 (
            .O(N__24985),
            .I(N__24982));
    LocalMux I__3485 (
            .O(N__24982),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__3484 (
            .O(N__24979),
            .I(N__24976));
    InMux I__3483 (
            .O(N__24976),
            .I(N__24973));
    LocalMux I__3482 (
            .O(N__24973),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__3481 (
            .O(N__24970),
            .I(N__24967));
    LocalMux I__3480 (
            .O(N__24967),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__3479 (
            .O(N__24964),
            .I(N__24961));
    InMux I__3478 (
            .O(N__24961),
            .I(N__24958));
    LocalMux I__3477 (
            .O(N__24958),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    InMux I__3476 (
            .O(N__24955),
            .I(N__24946));
    InMux I__3475 (
            .O(N__24954),
            .I(N__24946));
    InMux I__3474 (
            .O(N__24953),
            .I(N__24946));
    LocalMux I__3473 (
            .O(N__24946),
            .I(N__24943));
    Span4Mux_v I__3472 (
            .O(N__24943),
            .I(N__24939));
    InMux I__3471 (
            .O(N__24942),
            .I(N__24936));
    Span4Mux_v I__3470 (
            .O(N__24939),
            .I(N__24933));
    LocalMux I__3469 (
            .O(N__24936),
            .I(N__24930));
    Odrv4 I__3468 (
            .O(N__24933),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv12 I__3467 (
            .O(N__24930),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    CascadeMux I__3466 (
            .O(N__24925),
            .I(N__24922));
    InMux I__3465 (
            .O(N__24922),
            .I(N__24916));
    InMux I__3464 (
            .O(N__24921),
            .I(N__24916));
    LocalMux I__3463 (
            .O(N__24916),
            .I(N__24912));
    InMux I__3462 (
            .O(N__24915),
            .I(N__24909));
    Odrv4 I__3461 (
            .O(N__24912),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__3460 (
            .O(N__24909),
            .I(\current_shift_inst.un4_control_input1_29 ));
    CascadeMux I__3459 (
            .O(N__24904),
            .I(N__24901));
    InMux I__3458 (
            .O(N__24901),
            .I(N__24896));
    InMux I__3457 (
            .O(N__24900),
            .I(N__24891));
    InMux I__3456 (
            .O(N__24899),
            .I(N__24891));
    LocalMux I__3455 (
            .O(N__24896),
            .I(N__24888));
    LocalMux I__3454 (
            .O(N__24891),
            .I(N__24885));
    Span4Mux_v I__3453 (
            .O(N__24888),
            .I(N__24881));
    Span4Mux_h I__3452 (
            .O(N__24885),
            .I(N__24878));
    InMux I__3451 (
            .O(N__24884),
            .I(N__24875));
    Span4Mux_v I__3450 (
            .O(N__24881),
            .I(N__24872));
    Span4Mux_v I__3449 (
            .O(N__24878),
            .I(N__24869));
    LocalMux I__3448 (
            .O(N__24875),
            .I(N__24866));
    Odrv4 I__3447 (
            .O(N__24872),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__3446 (
            .O(N__24869),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv12 I__3445 (
            .O(N__24866),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    CascadeMux I__3444 (
            .O(N__24859),
            .I(N__24855));
    InMux I__3443 (
            .O(N__24858),
            .I(N__24851));
    InMux I__3442 (
            .O(N__24855),
            .I(N__24848));
    InMux I__3441 (
            .O(N__24854),
            .I(N__24845));
    LocalMux I__3440 (
            .O(N__24851),
            .I(\current_shift_inst.un4_control_input1_22 ));
    LocalMux I__3439 (
            .O(N__24848),
            .I(\current_shift_inst.un4_control_input1_22 ));
    LocalMux I__3438 (
            .O(N__24845),
            .I(\current_shift_inst.un4_control_input1_22 ));
    CascadeMux I__3437 (
            .O(N__24838),
            .I(N__24835));
    InMux I__3436 (
            .O(N__24835),
            .I(N__24830));
    InMux I__3435 (
            .O(N__24834),
            .I(N__24827));
    InMux I__3434 (
            .O(N__24833),
            .I(N__24824));
    LocalMux I__3433 (
            .O(N__24830),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__3432 (
            .O(N__24827),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__3431 (
            .O(N__24824),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__3430 (
            .O(N__24817),
            .I(N__24814));
    LocalMux I__3429 (
            .O(N__24814),
            .I(N__24809));
    InMux I__3428 (
            .O(N__24813),
            .I(N__24806));
    InMux I__3427 (
            .O(N__24812),
            .I(N__24803));
    Span4Mux_v I__3426 (
            .O(N__24809),
            .I(N__24795));
    LocalMux I__3425 (
            .O(N__24806),
            .I(N__24795));
    LocalMux I__3424 (
            .O(N__24803),
            .I(N__24795));
    InMux I__3423 (
            .O(N__24802),
            .I(N__24792));
    Odrv4 I__3422 (
            .O(N__24795),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__3421 (
            .O(N__24792),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    InMux I__3420 (
            .O(N__24787),
            .I(N__24783));
    CascadeMux I__3419 (
            .O(N__24786),
            .I(N__24779));
    LocalMux I__3418 (
            .O(N__24783),
            .I(N__24776));
    InMux I__3417 (
            .O(N__24782),
            .I(N__24771));
    InMux I__3416 (
            .O(N__24779),
            .I(N__24771));
    Span4Mux_v I__3415 (
            .O(N__24776),
            .I(N__24768));
    LocalMux I__3414 (
            .O(N__24771),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv4 I__3413 (
            .O(N__24768),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__3412 (
            .O(N__24763),
            .I(N__24757));
    InMux I__3411 (
            .O(N__24762),
            .I(N__24757));
    LocalMux I__3410 (
            .O(N__24757),
            .I(N__24753));
    InMux I__3409 (
            .O(N__24756),
            .I(N__24749));
    Sp12to4 I__3408 (
            .O(N__24753),
            .I(N__24746));
    InMux I__3407 (
            .O(N__24752),
            .I(N__24743));
    LocalMux I__3406 (
            .O(N__24749),
            .I(N__24740));
    Span12Mux_v I__3405 (
            .O(N__24746),
            .I(N__24737));
    LocalMux I__3404 (
            .O(N__24743),
            .I(N__24734));
    Span4Mux_v I__3403 (
            .O(N__24740),
            .I(N__24731));
    Odrv12 I__3402 (
            .O(N__24737),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__3401 (
            .O(N__24734),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__3400 (
            .O(N__24731),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    CascadeMux I__3399 (
            .O(N__24724),
            .I(N__24720));
    InMux I__3398 (
            .O(N__24723),
            .I(N__24715));
    InMux I__3397 (
            .O(N__24720),
            .I(N__24715));
    LocalMux I__3396 (
            .O(N__24715),
            .I(N__24712));
    Span4Mux_h I__3395 (
            .O(N__24712),
            .I(N__24708));
    InMux I__3394 (
            .O(N__24711),
            .I(N__24705));
    Span4Mux_v I__3393 (
            .O(N__24708),
            .I(N__24701));
    LocalMux I__3392 (
            .O(N__24705),
            .I(N__24698));
    InMux I__3391 (
            .O(N__24704),
            .I(N__24695));
    Odrv4 I__3390 (
            .O(N__24701),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__3389 (
            .O(N__24698),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__3388 (
            .O(N__24695),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    CascadeMux I__3387 (
            .O(N__24688),
            .I(N__24684));
    InMux I__3386 (
            .O(N__24687),
            .I(N__24680));
    InMux I__3385 (
            .O(N__24684),
            .I(N__24675));
    InMux I__3384 (
            .O(N__24683),
            .I(N__24675));
    LocalMux I__3383 (
            .O(N__24680),
            .I(N__24672));
    LocalMux I__3382 (
            .O(N__24675),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv12 I__3381 (
            .O(N__24672),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__3380 (
            .O(N__24667),
            .I(N__24664));
    LocalMux I__3379 (
            .O(N__24664),
            .I(N__24661));
    Odrv4 I__3378 (
            .O(N__24661),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__3377 (
            .O(N__24658),
            .I(N__24655));
    LocalMux I__3376 (
            .O(N__24655),
            .I(N__24652));
    Odrv4 I__3375 (
            .O(N__24652),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    InMux I__3374 (
            .O(N__24649),
            .I(N__24646));
    LocalMux I__3373 (
            .O(N__24646),
            .I(N__24643));
    Odrv4 I__3372 (
            .O(N__24643),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__3371 (
            .O(N__24640),
            .I(N__24637));
    LocalMux I__3370 (
            .O(N__24637),
            .I(N__24634));
    Odrv4 I__3369 (
            .O(N__24634),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__3368 (
            .O(N__24631),
            .I(N__24628));
    LocalMux I__3367 (
            .O(N__24628),
            .I(N__24625));
    Span4Mux_v I__3366 (
            .O(N__24625),
            .I(N__24622));
    Odrv4 I__3365 (
            .O(N__24622),
            .I(il_min_comp2_D1));
    InMux I__3364 (
            .O(N__24619),
            .I(N__24616));
    LocalMux I__3363 (
            .O(N__24616),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ));
    InMux I__3362 (
            .O(N__24613),
            .I(N__24610));
    LocalMux I__3361 (
            .O(N__24610),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__3360 (
            .O(N__24607),
            .I(N__24604));
    LocalMux I__3359 (
            .O(N__24604),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    InMux I__3358 (
            .O(N__24601),
            .I(N__24598));
    LocalMux I__3357 (
            .O(N__24598),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__3356 (
            .O(N__24595),
            .I(N__24592));
    LocalMux I__3355 (
            .O(N__24592),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    InMux I__3354 (
            .O(N__24589),
            .I(N__24586));
    LocalMux I__3353 (
            .O(N__24586),
            .I(N__24583));
    Span12Mux_h I__3352 (
            .O(N__24583),
            .I(N__24580));
    Odrv12 I__3351 (
            .O(N__24580),
            .I(il_max_comp1_c));
    CascadeMux I__3350 (
            .O(N__24577),
            .I(N__24574));
    InMux I__3349 (
            .O(N__24574),
            .I(N__24571));
    LocalMux I__3348 (
            .O(N__24571),
            .I(N__24566));
    InMux I__3347 (
            .O(N__24570),
            .I(N__24563));
    InMux I__3346 (
            .O(N__24569),
            .I(N__24560));
    Odrv4 I__3345 (
            .O(N__24566),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__3344 (
            .O(N__24563),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    LocalMux I__3343 (
            .O(N__24560),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ));
    InMux I__3342 (
            .O(N__24553),
            .I(N__24550));
    LocalMux I__3341 (
            .O(N__24550),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__3340 (
            .O(N__24547),
            .I(N__24544));
    LocalMux I__3339 (
            .O(N__24544),
            .I(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ));
    InMux I__3338 (
            .O(N__24541),
            .I(N__24538));
    LocalMux I__3337 (
            .O(N__24538),
            .I(\current_shift_inst.PI_CTRL.N_71 ));
    CascadeMux I__3336 (
            .O(N__24535),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ));
    CascadeMux I__3335 (
            .O(N__24532),
            .I(N__24529));
    InMux I__3334 (
            .O(N__24529),
            .I(N__24526));
    LocalMux I__3333 (
            .O(N__24526),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ));
    CascadeMux I__3332 (
            .O(N__24523),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10_cascade_ ));
    CascadeMux I__3331 (
            .O(N__24520),
            .I(N__24517));
    InMux I__3330 (
            .O(N__24517),
            .I(N__24514));
    LocalMux I__3329 (
            .O(N__24514),
            .I(N__24511));
    Odrv4 I__3328 (
            .O(N__24511),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    CascadeMux I__3327 (
            .O(N__24508),
            .I(N__24505));
    InMux I__3326 (
            .O(N__24505),
            .I(N__24500));
    InMux I__3325 (
            .O(N__24504),
            .I(N__24497));
    InMux I__3324 (
            .O(N__24503),
            .I(N__24494));
    LocalMux I__3323 (
            .O(N__24500),
            .I(N__24489));
    LocalMux I__3322 (
            .O(N__24497),
            .I(N__24489));
    LocalMux I__3321 (
            .O(N__24494),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__3320 (
            .O(N__24489),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__3319 (
            .O(N__24484),
            .I(bfn_8_24_0_));
    CascadeMux I__3318 (
            .O(N__24481),
            .I(N__24477));
    CascadeMux I__3317 (
            .O(N__24480),
            .I(N__24474));
    InMux I__3316 (
            .O(N__24477),
            .I(N__24470));
    InMux I__3315 (
            .O(N__24474),
            .I(N__24467));
    InMux I__3314 (
            .O(N__24473),
            .I(N__24464));
    LocalMux I__3313 (
            .O(N__24470),
            .I(N__24459));
    LocalMux I__3312 (
            .O(N__24467),
            .I(N__24459));
    LocalMux I__3311 (
            .O(N__24464),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__3310 (
            .O(N__24459),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__3309 (
            .O(N__24454),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__3308 (
            .O(N__24451),
            .I(N__24444));
    InMux I__3307 (
            .O(N__24450),
            .I(N__24444));
    InMux I__3306 (
            .O(N__24449),
            .I(N__24441));
    LocalMux I__3305 (
            .O(N__24444),
            .I(N__24438));
    LocalMux I__3304 (
            .O(N__24441),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__3303 (
            .O(N__24438),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__3302 (
            .O(N__24433),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    CascadeMux I__3301 (
            .O(N__24430),
            .I(N__24427));
    InMux I__3300 (
            .O(N__24427),
            .I(N__24422));
    InMux I__3299 (
            .O(N__24426),
            .I(N__24419));
    InMux I__3298 (
            .O(N__24425),
            .I(N__24416));
    LocalMux I__3297 (
            .O(N__24422),
            .I(N__24411));
    LocalMux I__3296 (
            .O(N__24419),
            .I(N__24411));
    LocalMux I__3295 (
            .O(N__24416),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__3294 (
            .O(N__24411),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__3293 (
            .O(N__24406),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    CascadeMux I__3292 (
            .O(N__24403),
            .I(N__24400));
    InMux I__3291 (
            .O(N__24400),
            .I(N__24396));
    InMux I__3290 (
            .O(N__24399),
            .I(N__24393));
    LocalMux I__3289 (
            .O(N__24396),
            .I(N__24390));
    LocalMux I__3288 (
            .O(N__24393),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__3287 (
            .O(N__24390),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__3286 (
            .O(N__24385),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__3285 (
            .O(N__24382),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__3284 (
            .O(N__24379),
            .I(N__24376));
    LocalMux I__3283 (
            .O(N__24376),
            .I(N__24372));
    InMux I__3282 (
            .O(N__24375),
            .I(N__24369));
    Span4Mux_h I__3281 (
            .O(N__24372),
            .I(N__24366));
    LocalMux I__3280 (
            .O(N__24369),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__3279 (
            .O(N__24366),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    InMux I__3278 (
            .O(N__24361),
            .I(N__24358));
    LocalMux I__3277 (
            .O(N__24358),
            .I(N__24355));
    Odrv12 I__3276 (
            .O(N__24355),
            .I(il_min_comp1_c));
    InMux I__3275 (
            .O(N__24352),
            .I(N__24345));
    InMux I__3274 (
            .O(N__24351),
            .I(N__24345));
    InMux I__3273 (
            .O(N__24350),
            .I(N__24342));
    LocalMux I__3272 (
            .O(N__24345),
            .I(N__24339));
    LocalMux I__3271 (
            .O(N__24342),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__3270 (
            .O(N__24339),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__3269 (
            .O(N__24334),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__3268 (
            .O(N__24331),
            .I(N__24328));
    InMux I__3267 (
            .O(N__24328),
            .I(N__24323));
    InMux I__3266 (
            .O(N__24327),
            .I(N__24320));
    InMux I__3265 (
            .O(N__24326),
            .I(N__24317));
    LocalMux I__3264 (
            .O(N__24323),
            .I(N__24312));
    LocalMux I__3263 (
            .O(N__24320),
            .I(N__24312));
    LocalMux I__3262 (
            .O(N__24317),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__3261 (
            .O(N__24312),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__3260 (
            .O(N__24307),
            .I(bfn_8_23_0_));
    CascadeMux I__3259 (
            .O(N__24304),
            .I(N__24300));
    CascadeMux I__3258 (
            .O(N__24303),
            .I(N__24297));
    InMux I__3257 (
            .O(N__24300),
            .I(N__24293));
    InMux I__3256 (
            .O(N__24297),
            .I(N__24290));
    InMux I__3255 (
            .O(N__24296),
            .I(N__24287));
    LocalMux I__3254 (
            .O(N__24293),
            .I(N__24282));
    LocalMux I__3253 (
            .O(N__24290),
            .I(N__24282));
    LocalMux I__3252 (
            .O(N__24287),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__3251 (
            .O(N__24282),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__3250 (
            .O(N__24277),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__3249 (
            .O(N__24274),
            .I(N__24267));
    InMux I__3248 (
            .O(N__24273),
            .I(N__24267));
    InMux I__3247 (
            .O(N__24272),
            .I(N__24264));
    LocalMux I__3246 (
            .O(N__24267),
            .I(N__24261));
    LocalMux I__3245 (
            .O(N__24264),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__3244 (
            .O(N__24261),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__3243 (
            .O(N__24256),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__3242 (
            .O(N__24253),
            .I(N__24250));
    InMux I__3241 (
            .O(N__24250),
            .I(N__24245));
    InMux I__3240 (
            .O(N__24249),
            .I(N__24242));
    InMux I__3239 (
            .O(N__24248),
            .I(N__24239));
    LocalMux I__3238 (
            .O(N__24245),
            .I(N__24234));
    LocalMux I__3237 (
            .O(N__24242),
            .I(N__24234));
    LocalMux I__3236 (
            .O(N__24239),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv4 I__3235 (
            .O(N__24234),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__3234 (
            .O(N__24229),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__3233 (
            .O(N__24226),
            .I(N__24222));
    InMux I__3232 (
            .O(N__24225),
            .I(N__24218));
    InMux I__3231 (
            .O(N__24222),
            .I(N__24215));
    InMux I__3230 (
            .O(N__24221),
            .I(N__24212));
    LocalMux I__3229 (
            .O(N__24218),
            .I(N__24207));
    LocalMux I__3228 (
            .O(N__24215),
            .I(N__24207));
    LocalMux I__3227 (
            .O(N__24212),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__3226 (
            .O(N__24207),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__3225 (
            .O(N__24202),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__3224 (
            .O(N__24199),
            .I(N__24196));
    InMux I__3223 (
            .O(N__24196),
            .I(N__24191));
    InMux I__3222 (
            .O(N__24195),
            .I(N__24188));
    InMux I__3221 (
            .O(N__24194),
            .I(N__24185));
    LocalMux I__3220 (
            .O(N__24191),
            .I(N__24180));
    LocalMux I__3219 (
            .O(N__24188),
            .I(N__24180));
    LocalMux I__3218 (
            .O(N__24185),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__3217 (
            .O(N__24180),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__3216 (
            .O(N__24175),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__3215 (
            .O(N__24172),
            .I(N__24168));
    CascadeMux I__3214 (
            .O(N__24171),
            .I(N__24165));
    InMux I__3213 (
            .O(N__24168),
            .I(N__24159));
    InMux I__3212 (
            .O(N__24165),
            .I(N__24159));
    InMux I__3211 (
            .O(N__24164),
            .I(N__24156));
    LocalMux I__3210 (
            .O(N__24159),
            .I(N__24153));
    LocalMux I__3209 (
            .O(N__24156),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__3208 (
            .O(N__24153),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__3207 (
            .O(N__24148),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__3206 (
            .O(N__24145),
            .I(N__24138));
    InMux I__3205 (
            .O(N__24144),
            .I(N__24138));
    InMux I__3204 (
            .O(N__24143),
            .I(N__24135));
    LocalMux I__3203 (
            .O(N__24138),
            .I(N__24132));
    LocalMux I__3202 (
            .O(N__24135),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__3201 (
            .O(N__24132),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__3200 (
            .O(N__24127),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__3199 (
            .O(N__24124),
            .I(N__24117));
    InMux I__3198 (
            .O(N__24123),
            .I(N__24117));
    InMux I__3197 (
            .O(N__24122),
            .I(N__24114));
    LocalMux I__3196 (
            .O(N__24117),
            .I(N__24111));
    LocalMux I__3195 (
            .O(N__24114),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__3194 (
            .O(N__24111),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__3193 (
            .O(N__24106),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__3192 (
            .O(N__24103),
            .I(N__24100));
    InMux I__3191 (
            .O(N__24100),
            .I(N__24095));
    InMux I__3190 (
            .O(N__24099),
            .I(N__24092));
    InMux I__3189 (
            .O(N__24098),
            .I(N__24089));
    LocalMux I__3188 (
            .O(N__24095),
            .I(N__24084));
    LocalMux I__3187 (
            .O(N__24092),
            .I(N__24084));
    LocalMux I__3186 (
            .O(N__24089),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv4 I__3185 (
            .O(N__24084),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__3184 (
            .O(N__24079),
            .I(bfn_8_22_0_));
    CascadeMux I__3183 (
            .O(N__24076),
            .I(N__24072));
    CascadeMux I__3182 (
            .O(N__24075),
            .I(N__24069));
    InMux I__3181 (
            .O(N__24072),
            .I(N__24066));
    InMux I__3180 (
            .O(N__24069),
            .I(N__24062));
    LocalMux I__3179 (
            .O(N__24066),
            .I(N__24059));
    InMux I__3178 (
            .O(N__24065),
            .I(N__24056));
    LocalMux I__3177 (
            .O(N__24062),
            .I(N__24051));
    Span4Mux_h I__3176 (
            .O(N__24059),
            .I(N__24051));
    LocalMux I__3175 (
            .O(N__24056),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__3174 (
            .O(N__24051),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__3173 (
            .O(N__24046),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__3172 (
            .O(N__24043),
            .I(N__24036));
    InMux I__3171 (
            .O(N__24042),
            .I(N__24036));
    InMux I__3170 (
            .O(N__24041),
            .I(N__24033));
    LocalMux I__3169 (
            .O(N__24036),
            .I(N__24030));
    LocalMux I__3168 (
            .O(N__24033),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__3167 (
            .O(N__24030),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__3166 (
            .O(N__24025),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    CascadeMux I__3165 (
            .O(N__24022),
            .I(N__24019));
    InMux I__3164 (
            .O(N__24019),
            .I(N__24014));
    InMux I__3163 (
            .O(N__24018),
            .I(N__24011));
    InMux I__3162 (
            .O(N__24017),
            .I(N__24008));
    LocalMux I__3161 (
            .O(N__24014),
            .I(N__24003));
    LocalMux I__3160 (
            .O(N__24011),
            .I(N__24003));
    LocalMux I__3159 (
            .O(N__24008),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__3158 (
            .O(N__24003),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__3157 (
            .O(N__23998),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__3156 (
            .O(N__23995),
            .I(N__23991));
    InMux I__3155 (
            .O(N__23994),
            .I(N__23987));
    InMux I__3154 (
            .O(N__23991),
            .I(N__23984));
    InMux I__3153 (
            .O(N__23990),
            .I(N__23981));
    LocalMux I__3152 (
            .O(N__23987),
            .I(N__23976));
    LocalMux I__3151 (
            .O(N__23984),
            .I(N__23976));
    LocalMux I__3150 (
            .O(N__23981),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__3149 (
            .O(N__23976),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__3148 (
            .O(N__23971),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__3147 (
            .O(N__23968),
            .I(N__23965));
    InMux I__3146 (
            .O(N__23965),
            .I(N__23960));
    InMux I__3145 (
            .O(N__23964),
            .I(N__23957));
    InMux I__3144 (
            .O(N__23963),
            .I(N__23954));
    LocalMux I__3143 (
            .O(N__23960),
            .I(N__23949));
    LocalMux I__3142 (
            .O(N__23957),
            .I(N__23949));
    LocalMux I__3141 (
            .O(N__23954),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__3140 (
            .O(N__23949),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__3139 (
            .O(N__23944),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__3138 (
            .O(N__23941),
            .I(N__23937));
    CascadeMux I__3137 (
            .O(N__23940),
            .I(N__23934));
    InMux I__3136 (
            .O(N__23937),
            .I(N__23928));
    InMux I__3135 (
            .O(N__23934),
            .I(N__23928));
    InMux I__3134 (
            .O(N__23933),
            .I(N__23925));
    LocalMux I__3133 (
            .O(N__23928),
            .I(N__23922));
    LocalMux I__3132 (
            .O(N__23925),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__3131 (
            .O(N__23922),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__3130 (
            .O(N__23917),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__3129 (
            .O(N__23914),
            .I(N__23909));
    InMux I__3128 (
            .O(N__23913),
            .I(N__23906));
    InMux I__3127 (
            .O(N__23912),
            .I(N__23903));
    LocalMux I__3126 (
            .O(N__23909),
            .I(N__23900));
    LocalMux I__3125 (
            .O(N__23906),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__3124 (
            .O(N__23903),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv4 I__3123 (
            .O(N__23900),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__3122 (
            .O(N__23893),
            .I(bfn_8_21_0_));
    InMux I__3121 (
            .O(N__23890),
            .I(N__23887));
    LocalMux I__3120 (
            .O(N__23887),
            .I(N__23882));
    InMux I__3119 (
            .O(N__23886),
            .I(N__23879));
    InMux I__3118 (
            .O(N__23885),
            .I(N__23876));
    Span4Mux_v I__3117 (
            .O(N__23882),
            .I(N__23871));
    LocalMux I__3116 (
            .O(N__23879),
            .I(N__23871));
    LocalMux I__3115 (
            .O(N__23876),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__3114 (
            .O(N__23871),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__3113 (
            .O(N__23866),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__3112 (
            .O(N__23863),
            .I(N__23859));
    CascadeMux I__3111 (
            .O(N__23862),
            .I(N__23856));
    InMux I__3110 (
            .O(N__23859),
            .I(N__23850));
    InMux I__3109 (
            .O(N__23856),
            .I(N__23850));
    InMux I__3108 (
            .O(N__23855),
            .I(N__23847));
    LocalMux I__3107 (
            .O(N__23850),
            .I(N__23844));
    LocalMux I__3106 (
            .O(N__23847),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv4 I__3105 (
            .O(N__23844),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__3104 (
            .O(N__23839),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    CascadeMux I__3103 (
            .O(N__23836),
            .I(N__23832));
    CascadeMux I__3102 (
            .O(N__23835),
            .I(N__23829));
    InMux I__3101 (
            .O(N__23832),
            .I(N__23823));
    InMux I__3100 (
            .O(N__23829),
            .I(N__23823));
    InMux I__3099 (
            .O(N__23828),
            .I(N__23820));
    LocalMux I__3098 (
            .O(N__23823),
            .I(N__23817));
    LocalMux I__3097 (
            .O(N__23820),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__3096 (
            .O(N__23817),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__3095 (
            .O(N__23812),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__3094 (
            .O(N__23809),
            .I(N__23806));
    InMux I__3093 (
            .O(N__23806),
            .I(N__23801));
    InMux I__3092 (
            .O(N__23805),
            .I(N__23798));
    InMux I__3091 (
            .O(N__23804),
            .I(N__23795));
    LocalMux I__3090 (
            .O(N__23801),
            .I(N__23790));
    LocalMux I__3089 (
            .O(N__23798),
            .I(N__23790));
    LocalMux I__3088 (
            .O(N__23795),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__3087 (
            .O(N__23790),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__3086 (
            .O(N__23785),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__3085 (
            .O(N__23782),
            .I(N__23779));
    InMux I__3084 (
            .O(N__23779),
            .I(N__23774));
    InMux I__3083 (
            .O(N__23778),
            .I(N__23771));
    InMux I__3082 (
            .O(N__23777),
            .I(N__23768));
    LocalMux I__3081 (
            .O(N__23774),
            .I(N__23763));
    LocalMux I__3080 (
            .O(N__23771),
            .I(N__23763));
    LocalMux I__3079 (
            .O(N__23768),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__3078 (
            .O(N__23763),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__3077 (
            .O(N__23758),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    CascadeMux I__3076 (
            .O(N__23755),
            .I(N__23752));
    InMux I__3075 (
            .O(N__23752),
            .I(N__23748));
    InMux I__3074 (
            .O(N__23751),
            .I(N__23745));
    LocalMux I__3073 (
            .O(N__23748),
            .I(N__23739));
    LocalMux I__3072 (
            .O(N__23745),
            .I(N__23739));
    InMux I__3071 (
            .O(N__23744),
            .I(N__23736));
    Span4Mux_h I__3070 (
            .O(N__23739),
            .I(N__23733));
    LocalMux I__3069 (
            .O(N__23736),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__3068 (
            .O(N__23733),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__3067 (
            .O(N__23728),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__3066 (
            .O(N__23725),
            .I(N__23722));
    LocalMux I__3065 (
            .O(N__23722),
            .I(N__23719));
    Span4Mux_v I__3064 (
            .O(N__23719),
            .I(N__23716));
    Odrv4 I__3063 (
            .O(N__23716),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__3062 (
            .O(N__23713),
            .I(N__23710));
    LocalMux I__3061 (
            .O(N__23710),
            .I(N__23707));
    Span4Mux_v I__3060 (
            .O(N__23707),
            .I(N__23704));
    Odrv4 I__3059 (
            .O(N__23704),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    CascadeMux I__3058 (
            .O(N__23701),
            .I(N__23698));
    InMux I__3057 (
            .O(N__23698),
            .I(N__23695));
    LocalMux I__3056 (
            .O(N__23695),
            .I(N__23692));
    Span4Mux_v I__3055 (
            .O(N__23692),
            .I(N__23689));
    Odrv4 I__3054 (
            .O(N__23689),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__3053 (
            .O(N__23686),
            .I(N__23683));
    LocalMux I__3052 (
            .O(N__23683),
            .I(N__23680));
    Odrv12 I__3051 (
            .O(N__23680),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__3050 (
            .O(N__23677),
            .I(N__23674));
    LocalMux I__3049 (
            .O(N__23674),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__3048 (
            .O(N__23671),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__3047 (
            .O(N__23668),
            .I(N__23665));
    LocalMux I__3046 (
            .O(N__23665),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__3045 (
            .O(N__23662),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__3044 (
            .O(N__23659),
            .I(N__23656));
    LocalMux I__3043 (
            .O(N__23656),
            .I(N__23653));
    Odrv4 I__3042 (
            .O(N__23653),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__3041 (
            .O(N__23650),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__3040 (
            .O(N__23647),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__3039 (
            .O(N__23644),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ));
    InMux I__3038 (
            .O(N__23641),
            .I(N__23638));
    LocalMux I__3037 (
            .O(N__23638),
            .I(N__23635));
    Odrv4 I__3036 (
            .O(N__23635),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__3035 (
            .O(N__23632),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__3034 (
            .O(N__23629),
            .I(N__23626));
    LocalMux I__3033 (
            .O(N__23626),
            .I(N__23623));
    Odrv4 I__3032 (
            .O(N__23623),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__3031 (
            .O(N__23620),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__3030 (
            .O(N__23617),
            .I(N__23614));
    LocalMux I__3029 (
            .O(N__23614),
            .I(N__23611));
    Odrv4 I__3028 (
            .O(N__23611),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__3027 (
            .O(N__23608),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__3026 (
            .O(N__23605),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__3025 (
            .O(N__23602),
            .I(N__23599));
    LocalMux I__3024 (
            .O(N__23599),
            .I(N__23596));
    Odrv4 I__3023 (
            .O(N__23596),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__3022 (
            .O(N__23593),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__3021 (
            .O(N__23590),
            .I(N__23587));
    LocalMux I__3020 (
            .O(N__23587),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__3019 (
            .O(N__23584),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__3018 (
            .O(N__23581),
            .I(N__23578));
    LocalMux I__3017 (
            .O(N__23578),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__3016 (
            .O(N__23575),
            .I(bfn_8_16_0_));
    InMux I__3015 (
            .O(N__23572),
            .I(N__23569));
    LocalMux I__3014 (
            .O(N__23569),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__3013 (
            .O(N__23566),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__3012 (
            .O(N__23563),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__3011 (
            .O(N__23560),
            .I(N__23557));
    LocalMux I__3010 (
            .O(N__23557),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__3009 (
            .O(N__23554),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__3008 (
            .O(N__23551),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__3007 (
            .O(N__23548),
            .I(N__23545));
    LocalMux I__3006 (
            .O(N__23545),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__3005 (
            .O(N__23542),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__3004 (
            .O(N__23539),
            .I(N__23536));
    LocalMux I__3003 (
            .O(N__23536),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__3002 (
            .O(N__23533),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__3001 (
            .O(N__23530),
            .I(N__23527));
    LocalMux I__3000 (
            .O(N__23527),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__2999 (
            .O(N__23524),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__2998 (
            .O(N__23521),
            .I(N__23518));
    LocalMux I__2997 (
            .O(N__23518),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__2996 (
            .O(N__23515),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__2995 (
            .O(N__23512),
            .I(N__23509));
    LocalMux I__2994 (
            .O(N__23509),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__2993 (
            .O(N__23506),
            .I(bfn_8_15_0_));
    InMux I__2992 (
            .O(N__23503),
            .I(N__23500));
    LocalMux I__2991 (
            .O(N__23500),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__2990 (
            .O(N__23497),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__2989 (
            .O(N__23494),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__2988 (
            .O(N__23491),
            .I(N__23488));
    LocalMux I__2987 (
            .O(N__23488),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__2986 (
            .O(N__23485),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__2985 (
            .O(N__23482),
            .I(N__23479));
    LocalMux I__2984 (
            .O(N__23479),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__2983 (
            .O(N__23476),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__2982 (
            .O(N__23473),
            .I(N__23470));
    LocalMux I__2981 (
            .O(N__23470),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__2980 (
            .O(N__23467),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__2979 (
            .O(N__23464),
            .I(N__23461));
    LocalMux I__2978 (
            .O(N__23461),
            .I(N__23458));
    Span4Mux_v I__2977 (
            .O(N__23458),
            .I(N__23455));
    Odrv4 I__2976 (
            .O(N__23455),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__2975 (
            .O(N__23452),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__2974 (
            .O(N__23449),
            .I(N__23446));
    LocalMux I__2973 (
            .O(N__23446),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__2972 (
            .O(N__23443),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__2971 (
            .O(N__23440),
            .I(N__23437));
    LocalMux I__2970 (
            .O(N__23437),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__2969 (
            .O(N__23434),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__2968 (
            .O(N__23431),
            .I(bfn_8_14_0_));
    CascadeMux I__2967 (
            .O(N__23428),
            .I(\current_shift_inst.PI_CTRL.N_72_cascade_ ));
    InMux I__2966 (
            .O(N__23425),
            .I(N__23422));
    LocalMux I__2965 (
            .O(N__23422),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    InMux I__2964 (
            .O(N__23419),
            .I(N__23416));
    LocalMux I__2963 (
            .O(N__23416),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__2962 (
            .O(N__23413),
            .I(N__23410));
    LocalMux I__2961 (
            .O(N__23410),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    InMux I__2960 (
            .O(N__23407),
            .I(N__23404));
    LocalMux I__2959 (
            .O(N__23404),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__2958 (
            .O(N__23401),
            .I(N__23398));
    LocalMux I__2957 (
            .O(N__23398),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__2956 (
            .O(N__23395),
            .I(N__23392));
    LocalMux I__2955 (
            .O(N__23392),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__2954 (
            .O(N__23389),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    InMux I__2953 (
            .O(N__23386),
            .I(N__23383));
    LocalMux I__2952 (
            .O(N__23383),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    InMux I__2951 (
            .O(N__23380),
            .I(N__23377));
    LocalMux I__2950 (
            .O(N__23377),
            .I(N__23374));
    Span12Mux_h I__2949 (
            .O(N__23374),
            .I(N__23371));
    Odrv12 I__2948 (
            .O(N__23371),
            .I(il_min_comp2_c));
    CascadeMux I__2947 (
            .O(N__23368),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ));
    InMux I__2946 (
            .O(N__23365),
            .I(N__23362));
    LocalMux I__2945 (
            .O(N__23362),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ));
    InMux I__2944 (
            .O(N__23359),
            .I(N__23356));
    LocalMux I__2943 (
            .O(N__23356),
            .I(N__23353));
    Span4Mux_h I__2942 (
            .O(N__23353),
            .I(N__23350));
    Odrv4 I__2941 (
            .O(N__23350),
            .I(il_max_comp2_D1));
    InMux I__2940 (
            .O(N__23347),
            .I(N__23344));
    LocalMux I__2939 (
            .O(N__23344),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    InMux I__2938 (
            .O(N__23341),
            .I(N__23338));
    LocalMux I__2937 (
            .O(N__23338),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    CascadeMux I__2936 (
            .O(N__23335),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_ ));
    CascadeMux I__2935 (
            .O(N__23332),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    InMux I__2934 (
            .O(N__23329),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__2933 (
            .O(N__23326),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__2932 (
            .O(N__23323),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__2931 (
            .O(N__23320),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__2930 (
            .O(N__23317),
            .I(bfn_7_22_0_));
    InMux I__2929 (
            .O(N__23314),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__2928 (
            .O(N__23311),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__2927 (
            .O(N__23308),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__2926 (
            .O(N__23305),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__2925 (
            .O(N__23302),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__2924 (
            .O(N__23299),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__2923 (
            .O(N__23296),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__2922 (
            .O(N__23293),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__2921 (
            .O(N__23290),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__2920 (
            .O(N__23287),
            .I(bfn_7_21_0_));
    InMux I__2919 (
            .O(N__23284),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__2918 (
            .O(N__23281),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__2917 (
            .O(N__23278),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__2916 (
            .O(N__23275),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__2915 (
            .O(N__23272),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__2914 (
            .O(N__23269),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__2913 (
            .O(N__23266),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    InMux I__2912 (
            .O(N__23263),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__2911 (
            .O(N__23260),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__2910 (
            .O(N__23257),
            .I(bfn_7_20_0_));
    InMux I__2909 (
            .O(N__23254),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__2908 (
            .O(N__23251),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__2907 (
            .O(N__23248),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__2906 (
            .O(N__23245),
            .I(N__23241));
    InMux I__2905 (
            .O(N__23244),
            .I(N__23238));
    LocalMux I__2904 (
            .O(N__23241),
            .I(N__23235));
    LocalMux I__2903 (
            .O(N__23238),
            .I(N__23232));
    Span4Mux_h I__2902 (
            .O(N__23235),
            .I(N__23227));
    Span4Mux_h I__2901 (
            .O(N__23232),
            .I(N__23227));
    Odrv4 I__2900 (
            .O(N__23227),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2899 (
            .O(N__23224),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    CascadeMux I__2898 (
            .O(N__23221),
            .I(N__23217));
    InMux I__2897 (
            .O(N__23220),
            .I(N__23214));
    InMux I__2896 (
            .O(N__23217),
            .I(N__23211));
    LocalMux I__2895 (
            .O(N__23214),
            .I(N__23206));
    LocalMux I__2894 (
            .O(N__23211),
            .I(N__23206));
    Span4Mux_h I__2893 (
            .O(N__23206),
            .I(N__23203));
    Span4Mux_h I__2892 (
            .O(N__23203),
            .I(N__23200));
    Odrv4 I__2891 (
            .O(N__23200),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2890 (
            .O(N__23197),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2889 (
            .O(N__23194),
            .I(N__23188));
    InMux I__2888 (
            .O(N__23193),
            .I(N__23188));
    LocalMux I__2887 (
            .O(N__23188),
            .I(N__23185));
    Odrv4 I__2886 (
            .O(N__23185),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2885 (
            .O(N__23182),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2884 (
            .O(N__23179),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2883 (
            .O(N__23176),
            .I(N__23172));
    InMux I__2882 (
            .O(N__23175),
            .I(N__23162));
    LocalMux I__2881 (
            .O(N__23172),
            .I(N__23159));
    InMux I__2880 (
            .O(N__23171),
            .I(N__23150));
    InMux I__2879 (
            .O(N__23170),
            .I(N__23150));
    InMux I__2878 (
            .O(N__23169),
            .I(N__23150));
    InMux I__2877 (
            .O(N__23168),
            .I(N__23150));
    InMux I__2876 (
            .O(N__23167),
            .I(N__23143));
    InMux I__2875 (
            .O(N__23166),
            .I(N__23143));
    InMux I__2874 (
            .O(N__23165),
            .I(N__23143));
    LocalMux I__2873 (
            .O(N__23162),
            .I(N__23139));
    Span4Mux_s3_h I__2872 (
            .O(N__23159),
            .I(N__23136));
    LocalMux I__2871 (
            .O(N__23150),
            .I(N__23133));
    LocalMux I__2870 (
            .O(N__23143),
            .I(N__23130));
    InMux I__2869 (
            .O(N__23142),
            .I(N__23127));
    Span4Mux_s3_h I__2868 (
            .O(N__23139),
            .I(N__23124));
    Span4Mux_v I__2867 (
            .O(N__23136),
            .I(N__23119));
    Span4Mux_s3_h I__2866 (
            .O(N__23133),
            .I(N__23119));
    Span4Mux_h I__2865 (
            .O(N__23130),
            .I(N__23114));
    LocalMux I__2864 (
            .O(N__23127),
            .I(N__23114));
    Span4Mux_h I__2863 (
            .O(N__23124),
            .I(N__23111));
    Span4Mux_h I__2862 (
            .O(N__23119),
            .I(N__23108));
    Span4Mux_h I__2861 (
            .O(N__23114),
            .I(N__23105));
    Odrv4 I__2860 (
            .O(N__23111),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2859 (
            .O(N__23108),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2858 (
            .O(N__23105),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__2857 (
            .O(N__23098),
            .I(N__23095));
    LocalMux I__2856 (
            .O(N__23095),
            .I(N__23091));
    InMux I__2855 (
            .O(N__23094),
            .I(N__23088));
    Span4Mux_v I__2854 (
            .O(N__23091),
            .I(N__23085));
    LocalMux I__2853 (
            .O(N__23088),
            .I(N__23082));
    Odrv4 I__2852 (
            .O(N__23085),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    Odrv12 I__2851 (
            .O(N__23082),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2850 (
            .O(N__23077),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__2849 (
            .O(N__23074),
            .I(N__23071));
    InMux I__2848 (
            .O(N__23071),
            .I(N__23067));
    InMux I__2847 (
            .O(N__23070),
            .I(N__23064));
    LocalMux I__2846 (
            .O(N__23067),
            .I(N__23059));
    LocalMux I__2845 (
            .O(N__23064),
            .I(N__23059));
    Odrv4 I__2844 (
            .O(N__23059),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2843 (
            .O(N__23056),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2842 (
            .O(N__23053),
            .I(N__23049));
    InMux I__2841 (
            .O(N__23052),
            .I(N__23046));
    LocalMux I__2840 (
            .O(N__23049),
            .I(N__23043));
    LocalMux I__2839 (
            .O(N__23046),
            .I(N__23040));
    Span4Mux_h I__2838 (
            .O(N__23043),
            .I(N__23037));
    Odrv4 I__2837 (
            .O(N__23040),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    Odrv4 I__2836 (
            .O(N__23037),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2835 (
            .O(N__23032),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2834 (
            .O(N__23029),
            .I(N__23023));
    InMux I__2833 (
            .O(N__23028),
            .I(N__23023));
    LocalMux I__2832 (
            .O(N__23023),
            .I(N__23020));
    Odrv4 I__2831 (
            .O(N__23020),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2830 (
            .O(N__23017),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2829 (
            .O(N__23014),
            .I(N__23008));
    InMux I__2828 (
            .O(N__23013),
            .I(N__23008));
    LocalMux I__2827 (
            .O(N__23008),
            .I(N__23005));
    Span4Mux_v I__2826 (
            .O(N__23005),
            .I(N__23002));
    Odrv4 I__2825 (
            .O(N__23002),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2824 (
            .O(N__22999),
            .I(bfn_7_12_0_));
    InMux I__2823 (
            .O(N__22996),
            .I(N__22990));
    InMux I__2822 (
            .O(N__22995),
            .I(N__22990));
    LocalMux I__2821 (
            .O(N__22990),
            .I(N__22987));
    Odrv4 I__2820 (
            .O(N__22987),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2819 (
            .O(N__22984),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ));
    CascadeMux I__2818 (
            .O(N__22981),
            .I(N__22977));
    CascadeMux I__2817 (
            .O(N__22980),
            .I(N__22974));
    InMux I__2816 (
            .O(N__22977),
            .I(N__22969));
    InMux I__2815 (
            .O(N__22974),
            .I(N__22969));
    LocalMux I__2814 (
            .O(N__22969),
            .I(N__22966));
    Odrv4 I__2813 (
            .O(N__22966),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2812 (
            .O(N__22963),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    CascadeMux I__2811 (
            .O(N__22960),
            .I(N__22956));
    InMux I__2810 (
            .O(N__22959),
            .I(N__22951));
    InMux I__2809 (
            .O(N__22956),
            .I(N__22951));
    LocalMux I__2808 (
            .O(N__22951),
            .I(N__22948));
    Odrv4 I__2807 (
            .O(N__22948),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2806 (
            .O(N__22945),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    CascadeMux I__2805 (
            .O(N__22942),
            .I(N__22938));
    InMux I__2804 (
            .O(N__22941),
            .I(N__22935));
    InMux I__2803 (
            .O(N__22938),
            .I(N__22932));
    LocalMux I__2802 (
            .O(N__22935),
            .I(N__22927));
    LocalMux I__2801 (
            .O(N__22932),
            .I(N__22927));
    Span4Mux_h I__2800 (
            .O(N__22927),
            .I(N__22924));
    Odrv4 I__2799 (
            .O(N__22924),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2798 (
            .O(N__22921),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2797 (
            .O(N__22918),
            .I(N__22914));
    InMux I__2796 (
            .O(N__22917),
            .I(N__22911));
    LocalMux I__2795 (
            .O(N__22914),
            .I(N__22906));
    LocalMux I__2794 (
            .O(N__22911),
            .I(N__22906));
    Span4Mux_v I__2793 (
            .O(N__22906),
            .I(N__22903));
    Odrv4 I__2792 (
            .O(N__22903),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2791 (
            .O(N__22900),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    CascadeMux I__2790 (
            .O(N__22897),
            .I(N__22893));
    CascadeMux I__2789 (
            .O(N__22896),
            .I(N__22890));
    InMux I__2788 (
            .O(N__22893),
            .I(N__22885));
    InMux I__2787 (
            .O(N__22890),
            .I(N__22885));
    LocalMux I__2786 (
            .O(N__22885),
            .I(N__22882));
    Span4Mux_v I__2785 (
            .O(N__22882),
            .I(N__22879));
    Odrv4 I__2784 (
            .O(N__22879),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2783 (
            .O(N__22876),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2782 (
            .O(N__22873),
            .I(N__22867));
    InMux I__2781 (
            .O(N__22872),
            .I(N__22867));
    LocalMux I__2780 (
            .O(N__22867),
            .I(N__22864));
    Span4Mux_h I__2779 (
            .O(N__22864),
            .I(N__22861));
    Odrv4 I__2778 (
            .O(N__22861),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2777 (
            .O(N__22858),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    CascadeMux I__2776 (
            .O(N__22855),
            .I(N__22852));
    InMux I__2775 (
            .O(N__22852),
            .I(N__22848));
    InMux I__2774 (
            .O(N__22851),
            .I(N__22845));
    LocalMux I__2773 (
            .O(N__22848),
            .I(N__22842));
    LocalMux I__2772 (
            .O(N__22845),
            .I(N__22839));
    Span4Mux_v I__2771 (
            .O(N__22842),
            .I(N__22836));
    Span4Mux_h I__2770 (
            .O(N__22839),
            .I(N__22833));
    Odrv4 I__2769 (
            .O(N__22836),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    Odrv4 I__2768 (
            .O(N__22833),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2767 (
            .O(N__22828),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__2766 (
            .O(N__22825),
            .I(N__22821));
    InMux I__2765 (
            .O(N__22824),
            .I(N__22818));
    LocalMux I__2764 (
            .O(N__22821),
            .I(N__22815));
    LocalMux I__2763 (
            .O(N__22818),
            .I(N__22812));
    Span4Mux_h I__2762 (
            .O(N__22815),
            .I(N__22809));
    Odrv4 I__2761 (
            .O(N__22812),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    Odrv4 I__2760 (
            .O(N__22809),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2759 (
            .O(N__22804),
            .I(bfn_7_11_0_));
    InMux I__2758 (
            .O(N__22801),
            .I(N__22797));
    InMux I__2757 (
            .O(N__22800),
            .I(N__22794));
    LocalMux I__2756 (
            .O(N__22797),
            .I(N__22791));
    LocalMux I__2755 (
            .O(N__22794),
            .I(N__22788));
    Span4Mux_h I__2754 (
            .O(N__22791),
            .I(N__22785));
    Odrv12 I__2753 (
            .O(N__22788),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    Odrv4 I__2752 (
            .O(N__22785),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2751 (
            .O(N__22780),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ));
    InMux I__2750 (
            .O(N__22777),
            .I(N__22773));
    InMux I__2749 (
            .O(N__22776),
            .I(N__22770));
    LocalMux I__2748 (
            .O(N__22773),
            .I(N__22767));
    LocalMux I__2747 (
            .O(N__22770),
            .I(N__22764));
    Span4Mux_h I__2746 (
            .O(N__22767),
            .I(N__22761));
    Span4Mux_h I__2745 (
            .O(N__22764),
            .I(N__22758));
    Odrv4 I__2744 (
            .O(N__22761),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    Odrv4 I__2743 (
            .O(N__22758),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2742 (
            .O(N__22753),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2741 (
            .O(N__22750),
            .I(N__22747));
    LocalMux I__2740 (
            .O(N__22747),
            .I(N__22743));
    InMux I__2739 (
            .O(N__22746),
            .I(N__22740));
    Span4Mux_h I__2738 (
            .O(N__22743),
            .I(N__22737));
    LocalMux I__2737 (
            .O(N__22740),
            .I(N__22734));
    Odrv4 I__2736 (
            .O(N__22737),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    Odrv4 I__2735 (
            .O(N__22734),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2734 (
            .O(N__22729),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2733 (
            .O(N__22726),
            .I(N__22721));
    InMux I__2732 (
            .O(N__22725),
            .I(N__22716));
    InMux I__2731 (
            .O(N__22724),
            .I(N__22716));
    LocalMux I__2730 (
            .O(N__22721),
            .I(N__22713));
    LocalMux I__2729 (
            .O(N__22716),
            .I(N__22710));
    Span4Mux_h I__2728 (
            .O(N__22713),
            .I(N__22707));
    Span4Mux_v I__2727 (
            .O(N__22710),
            .I(N__22704));
    Odrv4 I__2726 (
            .O(N__22707),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__2725 (
            .O(N__22704),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2724 (
            .O(N__22699),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__2723 (
            .O(N__22696),
            .I(N__22693));
    LocalMux I__2722 (
            .O(N__22693),
            .I(N__22687));
    InMux I__2721 (
            .O(N__22692),
            .I(N__22684));
    InMux I__2720 (
            .O(N__22691),
            .I(N__22679));
    InMux I__2719 (
            .O(N__22690),
            .I(N__22679));
    Span4Mux_v I__2718 (
            .O(N__22687),
            .I(N__22676));
    LocalMux I__2717 (
            .O(N__22684),
            .I(N__22671));
    LocalMux I__2716 (
            .O(N__22679),
            .I(N__22671));
    Span4Mux_h I__2715 (
            .O(N__22676),
            .I(N__22668));
    Span4Mux_h I__2714 (
            .O(N__22671),
            .I(N__22665));
    Odrv4 I__2713 (
            .O(N__22668),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2712 (
            .O(N__22665),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2711 (
            .O(N__22660),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    CascadeMux I__2710 (
            .O(N__22657),
            .I(N__22654));
    InMux I__2709 (
            .O(N__22654),
            .I(N__22651));
    LocalMux I__2708 (
            .O(N__22651),
            .I(N__22647));
    InMux I__2707 (
            .O(N__22650),
            .I(N__22644));
    Span4Mux_v I__2706 (
            .O(N__22647),
            .I(N__22641));
    LocalMux I__2705 (
            .O(N__22644),
            .I(N__22637));
    Span4Mux_s1_h I__2704 (
            .O(N__22641),
            .I(N__22634));
    InMux I__2703 (
            .O(N__22640),
            .I(N__22631));
    Span4Mux_v I__2702 (
            .O(N__22637),
            .I(N__22628));
    Span4Mux_h I__2701 (
            .O(N__22634),
            .I(N__22623));
    LocalMux I__2700 (
            .O(N__22631),
            .I(N__22623));
    Odrv4 I__2699 (
            .O(N__22628),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__2698 (
            .O(N__22623),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2697 (
            .O(N__22618),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2696 (
            .O(N__22615),
            .I(N__22612));
    LocalMux I__2695 (
            .O(N__22612),
            .I(N__22609));
    Span4Mux_s3_h I__2694 (
            .O(N__22609),
            .I(N__22604));
    InMux I__2693 (
            .O(N__22608),
            .I(N__22601));
    InMux I__2692 (
            .O(N__22607),
            .I(N__22598));
    Span4Mux_v I__2691 (
            .O(N__22604),
            .I(N__22593));
    LocalMux I__2690 (
            .O(N__22601),
            .I(N__22593));
    LocalMux I__2689 (
            .O(N__22598),
            .I(N__22590));
    Span4Mux_h I__2688 (
            .O(N__22593),
            .I(N__22587));
    Odrv4 I__2687 (
            .O(N__22590),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2686 (
            .O(N__22587),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2685 (
            .O(N__22582),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    CascadeMux I__2684 (
            .O(N__22579),
            .I(N__22575));
    CascadeMux I__2683 (
            .O(N__22578),
            .I(N__22572));
    InMux I__2682 (
            .O(N__22575),
            .I(N__22568));
    InMux I__2681 (
            .O(N__22572),
            .I(N__22565));
    InMux I__2680 (
            .O(N__22571),
            .I(N__22562));
    LocalMux I__2679 (
            .O(N__22568),
            .I(N__22559));
    LocalMux I__2678 (
            .O(N__22565),
            .I(N__22556));
    LocalMux I__2677 (
            .O(N__22562),
            .I(N__22551));
    Span4Mux_v I__2676 (
            .O(N__22559),
            .I(N__22551));
    Odrv12 I__2675 (
            .O(N__22556),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2674 (
            .O(N__22551),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2673 (
            .O(N__22546),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2672 (
            .O(N__22543),
            .I(N__22539));
    CascadeMux I__2671 (
            .O(N__22542),
            .I(N__22536));
    LocalMux I__2670 (
            .O(N__22539),
            .I(N__22533));
    InMux I__2669 (
            .O(N__22536),
            .I(N__22530));
    Span4Mux_h I__2668 (
            .O(N__22533),
            .I(N__22525));
    LocalMux I__2667 (
            .O(N__22530),
            .I(N__22525));
    Span4Mux_v I__2666 (
            .O(N__22525),
            .I(N__22521));
    InMux I__2665 (
            .O(N__22524),
            .I(N__22518));
    Sp12to4 I__2664 (
            .O(N__22521),
            .I(N__22513));
    LocalMux I__2663 (
            .O(N__22518),
            .I(N__22513));
    Odrv12 I__2662 (
            .O(N__22513),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2661 (
            .O(N__22510),
            .I(bfn_7_10_0_));
    CascadeMux I__2660 (
            .O(N__22507),
            .I(N__22504));
    InMux I__2659 (
            .O(N__22504),
            .I(N__22499));
    InMux I__2658 (
            .O(N__22503),
            .I(N__22496));
    InMux I__2657 (
            .O(N__22502),
            .I(N__22493));
    LocalMux I__2656 (
            .O(N__22499),
            .I(N__22490));
    LocalMux I__2655 (
            .O(N__22496),
            .I(N__22487));
    LocalMux I__2654 (
            .O(N__22493),
            .I(N__22484));
    Span4Mux_h I__2653 (
            .O(N__22490),
            .I(N__22479));
    Span4Mux_v I__2652 (
            .O(N__22487),
            .I(N__22479));
    Odrv12 I__2651 (
            .O(N__22484),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__2650 (
            .O(N__22479),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2649 (
            .O(N__22474),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ));
    InMux I__2648 (
            .O(N__22471),
            .I(N__22465));
    InMux I__2647 (
            .O(N__22470),
            .I(N__22465));
    LocalMux I__2646 (
            .O(N__22465),
            .I(N__22462));
    Span4Mux_h I__2645 (
            .O(N__22462),
            .I(N__22459));
    Odrv4 I__2644 (
            .O(N__22459),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2643 (
            .O(N__22456),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2642 (
            .O(N__22453),
            .I(N__22450));
    LocalMux I__2641 (
            .O(N__22450),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__2640 (
            .O(N__22447),
            .I(N__22444));
    LocalMux I__2639 (
            .O(N__22444),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ));
    InMux I__2638 (
            .O(N__22441),
            .I(N__22438));
    LocalMux I__2637 (
            .O(N__22438),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ));
    InMux I__2636 (
            .O(N__22435),
            .I(N__22432));
    LocalMux I__2635 (
            .O(N__22432),
            .I(N__22429));
    Span4Mux_s3_h I__2634 (
            .O(N__22429),
            .I(N__22426));
    Span4Mux_h I__2633 (
            .O(N__22426),
            .I(N__22423));
    Odrv4 I__2632 (
            .O(N__22423),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__2631 (
            .O(N__22420),
            .I(N__22417));
    LocalMux I__2630 (
            .O(N__22417),
            .I(N__22414));
    Span12Mux_s7_h I__2629 (
            .O(N__22414),
            .I(N__22411));
    Odrv12 I__2628 (
            .O(N__22411),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__2627 (
            .O(N__22408),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ));
    InMux I__2626 (
            .O(N__22405),
            .I(N__22402));
    LocalMux I__2625 (
            .O(N__22402),
            .I(N__22399));
    Span4Mux_h I__2624 (
            .O(N__22399),
            .I(N__22396));
    Odrv4 I__2623 (
            .O(N__22396),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2622 (
            .O(N__22393),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2621 (
            .O(N__22390),
            .I(N__22387));
    LocalMux I__2620 (
            .O(N__22387),
            .I(N__22384));
    Span4Mux_s1_h I__2619 (
            .O(N__22384),
            .I(N__22379));
    InMux I__2618 (
            .O(N__22383),
            .I(N__22376));
    InMux I__2617 (
            .O(N__22382),
            .I(N__22373));
    Span4Mux_h I__2616 (
            .O(N__22379),
            .I(N__22370));
    LocalMux I__2615 (
            .O(N__22376),
            .I(pwm_duty_input_3));
    LocalMux I__2614 (
            .O(N__22373),
            .I(pwm_duty_input_3));
    Odrv4 I__2613 (
            .O(N__22370),
            .I(pwm_duty_input_3));
    CascadeMux I__2612 (
            .O(N__22363),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ));
    CascadeMux I__2611 (
            .O(N__22360),
            .I(N__22352));
    CascadeMux I__2610 (
            .O(N__22359),
            .I(N__22349));
    InMux I__2609 (
            .O(N__22358),
            .I(N__22346));
    InMux I__2608 (
            .O(N__22357),
            .I(N__22335));
    InMux I__2607 (
            .O(N__22356),
            .I(N__22335));
    InMux I__2606 (
            .O(N__22355),
            .I(N__22335));
    InMux I__2605 (
            .O(N__22352),
            .I(N__22335));
    InMux I__2604 (
            .O(N__22349),
            .I(N__22335));
    LocalMux I__2603 (
            .O(N__22346),
            .I(N__22330));
    LocalMux I__2602 (
            .O(N__22335),
            .I(N__22330));
    Span4Mux_v I__2601 (
            .O(N__22330),
            .I(N__22326));
    InMux I__2600 (
            .O(N__22329),
            .I(N__22323));
    Span4Mux_h I__2599 (
            .O(N__22326),
            .I(N__22320));
    LocalMux I__2598 (
            .O(N__22323),
            .I(N__22317));
    Odrv4 I__2597 (
            .O(N__22320),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    Odrv4 I__2596 (
            .O(N__22317),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2595 (
            .O(N__22312),
            .I(N__22309));
    LocalMux I__2594 (
            .O(N__22309),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__2593 (
            .O(N__22306),
            .I(N__22303));
    LocalMux I__2592 (
            .O(N__22303),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__2591 (
            .O(N__22300),
            .I(N__22297));
    LocalMux I__2590 (
            .O(N__22297),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__2589 (
            .O(N__22294),
            .I(N__22291));
    LocalMux I__2588 (
            .O(N__22291),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ));
    InMux I__2587 (
            .O(N__22288),
            .I(N__22285));
    LocalMux I__2586 (
            .O(N__22285),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__2585 (
            .O(N__22282),
            .I(N__22279));
    LocalMux I__2584 (
            .O(N__22279),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__2583 (
            .O(N__22276),
            .I(N__22273));
    LocalMux I__2582 (
            .O(N__22273),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__2581 (
            .O(N__22270),
            .I(\current_shift_inst.PI_CTRL.N_53_cascade_ ));
    InMux I__2580 (
            .O(N__22267),
            .I(N__22261));
    InMux I__2579 (
            .O(N__22266),
            .I(N__22261));
    LocalMux I__2578 (
            .O(N__22261),
            .I(N__22258));
    Span4Mux_h I__2577 (
            .O(N__22258),
            .I(N__22254));
    InMux I__2576 (
            .O(N__22257),
            .I(N__22251));
    Odrv4 I__2575 (
            .O(N__22254),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    LocalMux I__2574 (
            .O(N__22251),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__2573 (
            .O(N__22246),
            .I(N__22243));
    LocalMux I__2572 (
            .O(N__22243),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    CascadeMux I__2571 (
            .O(N__22240),
            .I(N__22237));
    InMux I__2570 (
            .O(N__22237),
            .I(N__22234));
    LocalMux I__2569 (
            .O(N__22234),
            .I(\current_shift_inst.PI_CTRL.N_155 ));
    CascadeMux I__2568 (
            .O(N__22231),
            .I(N__22227));
    CascadeMux I__2567 (
            .O(N__22230),
            .I(N__22224));
    InMux I__2566 (
            .O(N__22227),
            .I(N__22218));
    InMux I__2565 (
            .O(N__22224),
            .I(N__22218));
    InMux I__2564 (
            .O(N__22223),
            .I(N__22215));
    LocalMux I__2563 (
            .O(N__22218),
            .I(N__22210));
    LocalMux I__2562 (
            .O(N__22215),
            .I(N__22210));
    Odrv4 I__2561 (
            .O(N__22210),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    ClkMux I__2560 (
            .O(N__22207),
            .I(N__22204));
    GlobalMux I__2559 (
            .O(N__22204),
            .I(N__22201));
    gio2CtrlBuf I__2558 (
            .O(N__22201),
            .I(delay_hc_input_c_g));
    InMux I__2557 (
            .O(N__22198),
            .I(N__22195));
    LocalMux I__2556 (
            .O(N__22195),
            .I(N__22192));
    Odrv12 I__2555 (
            .O(N__22192),
            .I(il_max_comp2_c));
    InMux I__2554 (
            .O(N__22189),
            .I(N__22186));
    LocalMux I__2553 (
            .O(N__22186),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ));
    CascadeMux I__2552 (
            .O(N__22183),
            .I(N__22179));
    CascadeMux I__2551 (
            .O(N__22182),
            .I(N__22176));
    InMux I__2550 (
            .O(N__22179),
            .I(N__22169));
    InMux I__2549 (
            .O(N__22176),
            .I(N__22169));
    InMux I__2548 (
            .O(N__22175),
            .I(N__22166));
    CascadeMux I__2547 (
            .O(N__22174),
            .I(N__22163));
    LocalMux I__2546 (
            .O(N__22169),
            .I(N__22160));
    LocalMux I__2545 (
            .O(N__22166),
            .I(N__22157));
    InMux I__2544 (
            .O(N__22163),
            .I(N__22153));
    Span4Mux_v I__2543 (
            .O(N__22160),
            .I(N__22148));
    Span4Mux_v I__2542 (
            .O(N__22157),
            .I(N__22148));
    InMux I__2541 (
            .O(N__22156),
            .I(N__22145));
    LocalMux I__2540 (
            .O(N__22153),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    Odrv4 I__2539 (
            .O(N__22148),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    LocalMux I__2538 (
            .O(N__22145),
            .I(\current_shift_inst.PI_CTRL.N_153 ));
    InMux I__2537 (
            .O(N__22138),
            .I(N__22134));
    InMux I__2536 (
            .O(N__22137),
            .I(N__22131));
    LocalMux I__2535 (
            .O(N__22134),
            .I(N__22128));
    LocalMux I__2534 (
            .O(N__22131),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    Odrv4 I__2533 (
            .O(N__22128),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    InMux I__2532 (
            .O(N__22123),
            .I(N__22115));
    InMux I__2531 (
            .O(N__22122),
            .I(N__22106));
    InMux I__2530 (
            .O(N__22121),
            .I(N__22106));
    InMux I__2529 (
            .O(N__22120),
            .I(N__22106));
    InMux I__2528 (
            .O(N__22119),
            .I(N__22106));
    CascadeMux I__2527 (
            .O(N__22118),
            .I(N__22103));
    LocalMux I__2526 (
            .O(N__22115),
            .I(N__22100));
    LocalMux I__2525 (
            .O(N__22106),
            .I(N__22097));
    InMux I__2524 (
            .O(N__22103),
            .I(N__22092));
    Span4Mux_v I__2523 (
            .O(N__22100),
            .I(N__22089));
    Span4Mux_h I__2522 (
            .O(N__22097),
            .I(N__22086));
    InMux I__2521 (
            .O(N__22096),
            .I(N__22081));
    InMux I__2520 (
            .O(N__22095),
            .I(N__22081));
    LocalMux I__2519 (
            .O(N__22092),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2518 (
            .O(N__22089),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    Odrv4 I__2517 (
            .O(N__22086),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    LocalMux I__2516 (
            .O(N__22081),
            .I(\current_shift_inst.PI_CTRL.N_53 ));
    InMux I__2515 (
            .O(N__22072),
            .I(N__22069));
    LocalMux I__2514 (
            .O(N__22069),
            .I(N__22066));
    Odrv4 I__2513 (
            .O(N__22066),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    InMux I__2512 (
            .O(N__22063),
            .I(N__22060));
    LocalMux I__2511 (
            .O(N__22060),
            .I(N__22055));
    InMux I__2510 (
            .O(N__22059),
            .I(N__22052));
    InMux I__2509 (
            .O(N__22058),
            .I(N__22049));
    Span4Mux_h I__2508 (
            .O(N__22055),
            .I(N__22046));
    LocalMux I__2507 (
            .O(N__22052),
            .I(N__22043));
    LocalMux I__2506 (
            .O(N__22049),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    Odrv4 I__2505 (
            .O(N__22046),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    Odrv4 I__2504 (
            .O(N__22043),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    CascadeMux I__2503 (
            .O(N__22036),
            .I(N__22033));
    InMux I__2502 (
            .O(N__22033),
            .I(N__22030));
    LocalMux I__2501 (
            .O(N__22030),
            .I(N__22027));
    Span4Mux_h I__2500 (
            .O(N__22027),
            .I(N__22023));
    InMux I__2499 (
            .O(N__22026),
            .I(N__22020));
    Odrv4 I__2498 (
            .O(N__22023),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    LocalMux I__2497 (
            .O(N__22020),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    CascadeMux I__2496 (
            .O(N__22015),
            .I(N__22010));
    CascadeMux I__2495 (
            .O(N__22014),
            .I(N__22006));
    CascadeMux I__2494 (
            .O(N__22013),
            .I(N__22000));
    InMux I__2493 (
            .O(N__22010),
            .I(N__21991));
    InMux I__2492 (
            .O(N__22009),
            .I(N__21991));
    InMux I__2491 (
            .O(N__22006),
            .I(N__21991));
    InMux I__2490 (
            .O(N__22005),
            .I(N__21988));
    CascadeMux I__2489 (
            .O(N__22004),
            .I(N__21985));
    CascadeMux I__2488 (
            .O(N__22003),
            .I(N__21982));
    InMux I__2487 (
            .O(N__22000),
            .I(N__21978));
    InMux I__2486 (
            .O(N__21999),
            .I(N__21975));
    InMux I__2485 (
            .O(N__21998),
            .I(N__21972));
    LocalMux I__2484 (
            .O(N__21991),
            .I(N__21969));
    LocalMux I__2483 (
            .O(N__21988),
            .I(N__21964));
    InMux I__2482 (
            .O(N__21985),
            .I(N__21961));
    InMux I__2481 (
            .O(N__21982),
            .I(N__21958));
    InMux I__2480 (
            .O(N__21981),
            .I(N__21955));
    LocalMux I__2479 (
            .O(N__21978),
            .I(N__21948));
    LocalMux I__2478 (
            .O(N__21975),
            .I(N__21948));
    LocalMux I__2477 (
            .O(N__21972),
            .I(N__21948));
    Span4Mux_v I__2476 (
            .O(N__21969),
            .I(N__21945));
    InMux I__2475 (
            .O(N__21968),
            .I(N__21940));
    InMux I__2474 (
            .O(N__21967),
            .I(N__21940));
    Span4Mux_h I__2473 (
            .O(N__21964),
            .I(N__21929));
    LocalMux I__2472 (
            .O(N__21961),
            .I(N__21929));
    LocalMux I__2471 (
            .O(N__21958),
            .I(N__21929));
    LocalMux I__2470 (
            .O(N__21955),
            .I(N__21929));
    Span4Mux_h I__2469 (
            .O(N__21948),
            .I(N__21929));
    Odrv4 I__2468 (
            .O(N__21945),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ));
    LocalMux I__2467 (
            .O(N__21940),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ));
    Odrv4 I__2466 (
            .O(N__21929),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ));
    InMux I__2465 (
            .O(N__21922),
            .I(N__21919));
    LocalMux I__2464 (
            .O(N__21919),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    InMux I__2463 (
            .O(N__21916),
            .I(N__21911));
    InMux I__2462 (
            .O(N__21915),
            .I(N__21908));
    InMux I__2461 (
            .O(N__21914),
            .I(N__21905));
    LocalMux I__2460 (
            .O(N__21911),
            .I(N__21902));
    LocalMux I__2459 (
            .O(N__21908),
            .I(N__21899));
    LocalMux I__2458 (
            .O(N__21905),
            .I(N__21896));
    Span4Mux_v I__2457 (
            .O(N__21902),
            .I(N__21893));
    Span4Mux_h I__2456 (
            .O(N__21899),
            .I(N__21890));
    Span4Mux_s1_h I__2455 (
            .O(N__21896),
            .I(N__21887));
    Odrv4 I__2454 (
            .O(N__21893),
            .I(pwm_duty_input_9));
    Odrv4 I__2453 (
            .O(N__21890),
            .I(pwm_duty_input_9));
    Odrv4 I__2452 (
            .O(N__21887),
            .I(pwm_duty_input_9));
    InMux I__2451 (
            .O(N__21880),
            .I(N__21875));
    CascadeMux I__2450 (
            .O(N__21879),
            .I(N__21872));
    InMux I__2449 (
            .O(N__21878),
            .I(N__21869));
    LocalMux I__2448 (
            .O(N__21875),
            .I(N__21866));
    InMux I__2447 (
            .O(N__21872),
            .I(N__21863));
    LocalMux I__2446 (
            .O(N__21869),
            .I(N__21860));
    Span4Mux_h I__2445 (
            .O(N__21866),
            .I(N__21857));
    LocalMux I__2444 (
            .O(N__21863),
            .I(N__21854));
    Span4Mux_s2_h I__2443 (
            .O(N__21860),
            .I(N__21851));
    Odrv4 I__2442 (
            .O(N__21857),
            .I(pwm_duty_input_6));
    Odrv4 I__2441 (
            .O(N__21854),
            .I(pwm_duty_input_6));
    Odrv4 I__2440 (
            .O(N__21851),
            .I(pwm_duty_input_6));
    InMux I__2439 (
            .O(N__21844),
            .I(N__21841));
    LocalMux I__2438 (
            .O(N__21841),
            .I(N__21836));
    InMux I__2437 (
            .O(N__21840),
            .I(N__21833));
    InMux I__2436 (
            .O(N__21839),
            .I(N__21830));
    Span4Mux_v I__2435 (
            .O(N__21836),
            .I(N__21825));
    LocalMux I__2434 (
            .O(N__21833),
            .I(N__21825));
    LocalMux I__2433 (
            .O(N__21830),
            .I(N__21822));
    Odrv4 I__2432 (
            .O(N__21825),
            .I(pwm_duty_input_8));
    Odrv4 I__2431 (
            .O(N__21822),
            .I(pwm_duty_input_8));
    CascadeMux I__2430 (
            .O(N__21817),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ));
    InMux I__2429 (
            .O(N__21814),
            .I(N__21808));
    InMux I__2428 (
            .O(N__21813),
            .I(N__21808));
    LocalMux I__2427 (
            .O(N__21808),
            .I(N__21797));
    InMux I__2426 (
            .O(N__21807),
            .I(N__21794));
    InMux I__2425 (
            .O(N__21806),
            .I(N__21779));
    InMux I__2424 (
            .O(N__21805),
            .I(N__21779));
    InMux I__2423 (
            .O(N__21804),
            .I(N__21779));
    InMux I__2422 (
            .O(N__21803),
            .I(N__21779));
    InMux I__2421 (
            .O(N__21802),
            .I(N__21779));
    InMux I__2420 (
            .O(N__21801),
            .I(N__21779));
    InMux I__2419 (
            .O(N__21800),
            .I(N__21779));
    Span4Mux_h I__2418 (
            .O(N__21797),
            .I(N__21774));
    LocalMux I__2417 (
            .O(N__21794),
            .I(N__21774));
    LocalMux I__2416 (
            .O(N__21779),
            .I(\pwm_generator_inst.N_17 ));
    Odrv4 I__2415 (
            .O(N__21774),
            .I(\pwm_generator_inst.N_17 ));
    InMux I__2414 (
            .O(N__21769),
            .I(N__21765));
    InMux I__2413 (
            .O(N__21768),
            .I(N__21762));
    LocalMux I__2412 (
            .O(N__21765),
            .I(N__21756));
    LocalMux I__2411 (
            .O(N__21762),
            .I(N__21756));
    InMux I__2410 (
            .O(N__21761),
            .I(N__21753));
    Span4Mux_s3_h I__2409 (
            .O(N__21756),
            .I(N__21750));
    LocalMux I__2408 (
            .O(N__21753),
            .I(\current_shift_inst.PI_CTRL.N_154 ));
    Odrv4 I__2407 (
            .O(N__21750),
            .I(\current_shift_inst.PI_CTRL.N_154 ));
    InMux I__2406 (
            .O(N__21745),
            .I(N__21741));
    InMux I__2405 (
            .O(N__21744),
            .I(N__21738));
    LocalMux I__2404 (
            .O(N__21741),
            .I(N__21735));
    LocalMux I__2403 (
            .O(N__21738),
            .I(N__21730));
    Span4Mux_v I__2402 (
            .O(N__21735),
            .I(N__21730));
    Odrv4 I__2401 (
            .O(N__21730),
            .I(pwm_duty_input_2));
    CascadeMux I__2400 (
            .O(N__21727),
            .I(N__21724));
    InMux I__2399 (
            .O(N__21724),
            .I(N__21719));
    InMux I__2398 (
            .O(N__21723),
            .I(N__21716));
    InMux I__2397 (
            .O(N__21722),
            .I(N__21713));
    LocalMux I__2396 (
            .O(N__21719),
            .I(N__21710));
    LocalMux I__2395 (
            .O(N__21716),
            .I(N__21707));
    LocalMux I__2394 (
            .O(N__21713),
            .I(N__21704));
    Sp12to4 I__2393 (
            .O(N__21710),
            .I(N__21699));
    Span12Mux_v I__2392 (
            .O(N__21707),
            .I(N__21699));
    Span4Mux_s1_h I__2391 (
            .O(N__21704),
            .I(N__21696));
    Odrv12 I__2390 (
            .O(N__21699),
            .I(pwm_duty_input_7));
    Odrv4 I__2389 (
            .O(N__21696),
            .I(pwm_duty_input_7));
    InMux I__2388 (
            .O(N__21691),
            .I(N__21687));
    InMux I__2387 (
            .O(N__21690),
            .I(N__21683));
    LocalMux I__2386 (
            .O(N__21687),
            .I(N__21680));
    InMux I__2385 (
            .O(N__21686),
            .I(N__21677));
    LocalMux I__2384 (
            .O(N__21683),
            .I(N__21674));
    Span4Mux_v I__2383 (
            .O(N__21680),
            .I(N__21669));
    LocalMux I__2382 (
            .O(N__21677),
            .I(N__21669));
    Span4Mux_s1_h I__2381 (
            .O(N__21674),
            .I(N__21666));
    Odrv4 I__2380 (
            .O(N__21669),
            .I(pwm_duty_input_5));
    Odrv4 I__2379 (
            .O(N__21666),
            .I(pwm_duty_input_5));
    InMux I__2378 (
            .O(N__21661),
            .I(N__21658));
    LocalMux I__2377 (
            .O(N__21658),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ));
    InMux I__2376 (
            .O(N__21655),
            .I(N__21652));
    LocalMux I__2375 (
            .O(N__21652),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    CascadeMux I__2374 (
            .O(N__21649),
            .I(N__21645));
    InMux I__2373 (
            .O(N__21648),
            .I(N__21641));
    InMux I__2372 (
            .O(N__21645),
            .I(N__21638));
    InMux I__2371 (
            .O(N__21644),
            .I(N__21635));
    LocalMux I__2370 (
            .O(N__21641),
            .I(N__21632));
    LocalMux I__2369 (
            .O(N__21638),
            .I(N__21629));
    LocalMux I__2368 (
            .O(N__21635),
            .I(N__21626));
    Span4Mux_v I__2367 (
            .O(N__21632),
            .I(N__21619));
    Span4Mux_h I__2366 (
            .O(N__21629),
            .I(N__21619));
    Span4Mux_v I__2365 (
            .O(N__21626),
            .I(N__21619));
    Odrv4 I__2364 (
            .O(N__21619),
            .I(pwm_duty_input_4));
    InMux I__2363 (
            .O(N__21616),
            .I(N__21613));
    LocalMux I__2362 (
            .O(N__21613),
            .I(N__21610));
    Odrv4 I__2361 (
            .O(N__21610),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__2360 (
            .O(N__21607),
            .I(N__21583));
    InMux I__2359 (
            .O(N__21606),
            .I(N__21583));
    InMux I__2358 (
            .O(N__21605),
            .I(N__21583));
    InMux I__2357 (
            .O(N__21604),
            .I(N__21583));
    InMux I__2356 (
            .O(N__21603),
            .I(N__21583));
    InMux I__2355 (
            .O(N__21602),
            .I(N__21583));
    InMux I__2354 (
            .O(N__21601),
            .I(N__21583));
    InMux I__2353 (
            .O(N__21600),
            .I(N__21580));
    InMux I__2352 (
            .O(N__21599),
            .I(N__21575));
    InMux I__2351 (
            .O(N__21598),
            .I(N__21575));
    LocalMux I__2350 (
            .O(N__21583),
            .I(N__21568));
    LocalMux I__2349 (
            .O(N__21580),
            .I(N__21568));
    LocalMux I__2348 (
            .O(N__21575),
            .I(N__21568));
    Span4Mux_v I__2347 (
            .O(N__21568),
            .I(N__21565));
    Odrv4 I__2346 (
            .O(N__21565),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__2345 (
            .O(N__21562),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ));
    CascadeMux I__2344 (
            .O(N__21559),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ));
    CascadeMux I__2343 (
            .O(N__21556),
            .I(N__21553));
    InMux I__2342 (
            .O(N__21553),
            .I(N__21550));
    LocalMux I__2341 (
            .O(N__21550),
            .I(N__21547));
    Odrv4 I__2340 (
            .O(N__21547),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671 ));
    CascadeMux I__2339 (
            .O(N__21544),
            .I(N__21541));
    InMux I__2338 (
            .O(N__21541),
            .I(N__21538));
    LocalMux I__2337 (
            .O(N__21538),
            .I(N__21535));
    Odrv4 I__2336 (
            .O(N__21535),
            .I(\pwm_generator_inst.threshold_9 ));
    CascadeMux I__2335 (
            .O(N__21532),
            .I(N__21529));
    InMux I__2334 (
            .O(N__21529),
            .I(N__21526));
    LocalMux I__2333 (
            .O(N__21526),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1 ));
    CascadeMux I__2332 (
            .O(N__21523),
            .I(N__21520));
    InMux I__2331 (
            .O(N__21520),
            .I(N__21517));
    LocalMux I__2330 (
            .O(N__21517),
            .I(\pwm_generator_inst.threshold_5 ));
    InMux I__2329 (
            .O(N__21514),
            .I(N__21511));
    LocalMux I__2328 (
            .O(N__21511),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61 ));
    CascadeMux I__2327 (
            .O(N__21508),
            .I(N__21505));
    InMux I__2326 (
            .O(N__21505),
            .I(N__21502));
    LocalMux I__2325 (
            .O(N__21502),
            .I(N__21499));
    Odrv4 I__2324 (
            .O(N__21499),
            .I(\pwm_generator_inst.un14_counter_6 ));
    CascadeMux I__2323 (
            .O(N__21496),
            .I(N__21493));
    InMux I__2322 (
            .O(N__21493),
            .I(N__21490));
    LocalMux I__2321 (
            .O(N__21490),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1 ));
    CascadeMux I__2320 (
            .O(N__21487),
            .I(N__21484));
    InMux I__2319 (
            .O(N__21484),
            .I(N__21481));
    LocalMux I__2318 (
            .O(N__21481),
            .I(\pwm_generator_inst.threshold_4 ));
    InMux I__2317 (
            .O(N__21478),
            .I(N__21475));
    LocalMux I__2316 (
            .O(N__21475),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791 ));
    CascadeMux I__2315 (
            .O(N__21472),
            .I(N__21469));
    InMux I__2314 (
            .O(N__21469),
            .I(N__21466));
    LocalMux I__2313 (
            .O(N__21466),
            .I(\pwm_generator_inst.un14_counter_1 ));
    CascadeMux I__2312 (
            .O(N__21463),
            .I(N__21460));
    InMux I__2311 (
            .O(N__21460),
            .I(N__21457));
    LocalMux I__2310 (
            .O(N__21457),
            .I(N__21454));
    Span4Mux_h I__2309 (
            .O(N__21454),
            .I(N__21451));
    Odrv4 I__2308 (
            .O(N__21451),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271 ));
    CascadeMux I__2307 (
            .O(N__21448),
            .I(N__21445));
    InMux I__2306 (
            .O(N__21445),
            .I(N__21442));
    LocalMux I__2305 (
            .O(N__21442),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__2304 (
            .O(N__21439),
            .I(N__21436));
    LocalMux I__2303 (
            .O(N__21436),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61 ));
    CascadeMux I__2302 (
            .O(N__21433),
            .I(N__21425));
    CascadeMux I__2301 (
            .O(N__21432),
            .I(N__21420));
    CascadeMux I__2300 (
            .O(N__21431),
            .I(N__21415));
    CascadeMux I__2299 (
            .O(N__21430),
            .I(N__21412));
    CascadeMux I__2298 (
            .O(N__21429),
            .I(N__21403));
    CascadeMux I__2297 (
            .O(N__21428),
            .I(N__21400));
    InMux I__2296 (
            .O(N__21425),
            .I(N__21397));
    InMux I__2295 (
            .O(N__21424),
            .I(N__21382));
    InMux I__2294 (
            .O(N__21423),
            .I(N__21382));
    InMux I__2293 (
            .O(N__21420),
            .I(N__21382));
    InMux I__2292 (
            .O(N__21419),
            .I(N__21382));
    InMux I__2291 (
            .O(N__21418),
            .I(N__21382));
    InMux I__2290 (
            .O(N__21415),
            .I(N__21382));
    InMux I__2289 (
            .O(N__21412),
            .I(N__21382));
    InMux I__2288 (
            .O(N__21411),
            .I(N__21379));
    InMux I__2287 (
            .O(N__21410),
            .I(N__21373));
    InMux I__2286 (
            .O(N__21409),
            .I(N__21373));
    InMux I__2285 (
            .O(N__21408),
            .I(N__21366));
    InMux I__2284 (
            .O(N__21407),
            .I(N__21366));
    InMux I__2283 (
            .O(N__21406),
            .I(N__21366));
    InMux I__2282 (
            .O(N__21403),
            .I(N__21361));
    InMux I__2281 (
            .O(N__21400),
            .I(N__21361));
    LocalMux I__2280 (
            .O(N__21397),
            .I(N__21356));
    LocalMux I__2279 (
            .O(N__21382),
            .I(N__21356));
    LocalMux I__2278 (
            .O(N__21379),
            .I(N__21338));
    InMux I__2277 (
            .O(N__21378),
            .I(N__21335));
    LocalMux I__2276 (
            .O(N__21373),
            .I(N__21330));
    LocalMux I__2275 (
            .O(N__21366),
            .I(N__21330));
    LocalMux I__2274 (
            .O(N__21361),
            .I(N__21325));
    Span4Mux_v I__2273 (
            .O(N__21356),
            .I(N__21325));
    InMux I__2272 (
            .O(N__21355),
            .I(N__21308));
    InMux I__2271 (
            .O(N__21354),
            .I(N__21308));
    InMux I__2270 (
            .O(N__21353),
            .I(N__21308));
    InMux I__2269 (
            .O(N__21352),
            .I(N__21308));
    InMux I__2268 (
            .O(N__21351),
            .I(N__21308));
    InMux I__2267 (
            .O(N__21350),
            .I(N__21308));
    InMux I__2266 (
            .O(N__21349),
            .I(N__21308));
    InMux I__2265 (
            .O(N__21348),
            .I(N__21308));
    InMux I__2264 (
            .O(N__21347),
            .I(N__21293));
    InMux I__2263 (
            .O(N__21346),
            .I(N__21293));
    InMux I__2262 (
            .O(N__21345),
            .I(N__21293));
    InMux I__2261 (
            .O(N__21344),
            .I(N__21293));
    InMux I__2260 (
            .O(N__21343),
            .I(N__21293));
    InMux I__2259 (
            .O(N__21342),
            .I(N__21293));
    InMux I__2258 (
            .O(N__21341),
            .I(N__21293));
    Span12Mux_v I__2257 (
            .O(N__21338),
            .I(N__21286));
    LocalMux I__2256 (
            .O(N__21335),
            .I(N__21286));
    Span12Mux_s1_h I__2255 (
            .O(N__21330),
            .I(N__21286));
    Odrv4 I__2254 (
            .O(N__21325),
            .I(N_19_1));
    LocalMux I__2253 (
            .O(N__21308),
            .I(N_19_1));
    LocalMux I__2252 (
            .O(N__21293),
            .I(N_19_1));
    Odrv12 I__2251 (
            .O(N__21286),
            .I(N_19_1));
    InMux I__2250 (
            .O(N__21277),
            .I(N__21274));
    LocalMux I__2249 (
            .O(N__21274),
            .I(\pwm_generator_inst.un14_counter_7 ));
    InMux I__2248 (
            .O(N__21271),
            .I(N__21268));
    LocalMux I__2247 (
            .O(N__21268),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ));
    InMux I__2246 (
            .O(N__21265),
            .I(N__21262));
    LocalMux I__2245 (
            .O(N__21262),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    InMux I__2244 (
            .O(N__21259),
            .I(N__21256));
    LocalMux I__2243 (
            .O(N__21256),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    InMux I__2242 (
            .O(N__21253),
            .I(N__21250));
    LocalMux I__2241 (
            .O(N__21250),
            .I(N__21247));
    Span4Mux_s2_h I__2240 (
            .O(N__21247),
            .I(N__21243));
    InMux I__2239 (
            .O(N__21246),
            .I(N__21240));
    Odrv4 I__2238 (
            .O(N__21243),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__2237 (
            .O(N__21240),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__2236 (
            .O(N__21235),
            .I(N__21232));
    InMux I__2235 (
            .O(N__21232),
            .I(N__21229));
    LocalMux I__2234 (
            .O(N__21229),
            .I(N__21226));
    Span4Mux_v I__2233 (
            .O(N__21226),
            .I(N__21223));
    Odrv4 I__2232 (
            .O(N__21223),
            .I(\current_shift_inst.PI_CTRL.N_149 ));
    InMux I__2231 (
            .O(N__21220),
            .I(N__21217));
    LocalMux I__2230 (
            .O(N__21217),
            .I(N__21213));
    InMux I__2229 (
            .O(N__21216),
            .I(N__21210));
    Odrv4 I__2228 (
            .O(N__21213),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    LocalMux I__2227 (
            .O(N__21210),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    InMux I__2226 (
            .O(N__21205),
            .I(N__21201));
    InMux I__2225 (
            .O(N__21204),
            .I(N__21198));
    LocalMux I__2224 (
            .O(N__21201),
            .I(N__21192));
    LocalMux I__2223 (
            .O(N__21198),
            .I(N__21192));
    InMux I__2222 (
            .O(N__21197),
            .I(N__21189));
    Span4Mux_v I__2221 (
            .O(N__21192),
            .I(N__21186));
    LocalMux I__2220 (
            .O(N__21189),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__2219 (
            .O(N__21186),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__2218 (
            .O(N__21181),
            .I(N__21178));
    LocalMux I__2217 (
            .O(N__21178),
            .I(N__21175));
    Glb2LocalMux I__2216 (
            .O(N__21175),
            .I(N__21172));
    GlobalMux I__2215 (
            .O(N__21172),
            .I(clk_12mhz));
    IoInMux I__2214 (
            .O(N__21169),
            .I(N__21166));
    LocalMux I__2213 (
            .O(N__21166),
            .I(N__21163));
    Span4Mux_s0_v I__2212 (
            .O(N__21163),
            .I(N__21160));
    Span4Mux_h I__2211 (
            .O(N__21160),
            .I(N__21157));
    Odrv4 I__2210 (
            .O(N__21157),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2209 (
            .O(N__21154),
            .I(N__21151));
    LocalMux I__2208 (
            .O(N__21151),
            .I(N__21148));
    Odrv4 I__2207 (
            .O(N__21148),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31 ));
    CascadeMux I__2206 (
            .O(N__21145),
            .I(N__21142));
    InMux I__2205 (
            .O(N__21142),
            .I(N__21139));
    LocalMux I__2204 (
            .O(N__21139),
            .I(\pwm_generator_inst.threshold_0 ));
    InMux I__2203 (
            .O(N__21136),
            .I(N__21133));
    LocalMux I__2202 (
            .O(N__21133),
            .I(N__21130));
    Span4Mux_h I__2201 (
            .O(N__21130),
            .I(N__21127));
    Odrv4 I__2200 (
            .O(N__21127),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__2199 (
            .O(N__21124),
            .I(N__21121));
    LocalMux I__2198 (
            .O(N__21121),
            .I(N__21118));
    Odrv4 I__2197 (
            .O(N__21118),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1 ));
    InMux I__2196 (
            .O(N__21115),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__2195 (
            .O(N__21112),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    InMux I__2194 (
            .O(N__21109),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__2193 (
            .O(N__21106),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__2192 (
            .O(N__21103),
            .I(N__21100));
    LocalMux I__2191 (
            .O(N__21100),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    InMux I__2190 (
            .O(N__21097),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    InMux I__2189 (
            .O(N__21094),
            .I(N__21091));
    LocalMux I__2188 (
            .O(N__21091),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__2187 (
            .O(N__21088),
            .I(bfn_3_10_0_));
    InMux I__2186 (
            .O(N__21085),
            .I(N__21082));
    LocalMux I__2185 (
            .O(N__21082),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    InMux I__2184 (
            .O(N__21079),
            .I(N__21076));
    LocalMux I__2183 (
            .O(N__21076),
            .I(N__21073));
    Span4Mux_h I__2182 (
            .O(N__21073),
            .I(N__21070));
    Odrv4 I__2181 (
            .O(N__21070),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8 ));
    InMux I__2180 (
            .O(N__21067),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    InMux I__2179 (
            .O(N__21064),
            .I(N__21060));
    InMux I__2178 (
            .O(N__21063),
            .I(N__21057));
    LocalMux I__2177 (
            .O(N__21060),
            .I(N__21054));
    LocalMux I__2176 (
            .O(N__21057),
            .I(N__21051));
    Odrv4 I__2175 (
            .O(N__21054),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8 ));
    Odrv4 I__2174 (
            .O(N__21051),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8 ));
    CascadeMux I__2173 (
            .O(N__21046),
            .I(N__21042));
    InMux I__2172 (
            .O(N__21045),
            .I(N__21038));
    InMux I__2171 (
            .O(N__21042),
            .I(N__21035));
    InMux I__2170 (
            .O(N__21041),
            .I(N__21032));
    LocalMux I__2169 (
            .O(N__21038),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__2168 (
            .O(N__21035),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__2167 (
            .O(N__21032),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    InMux I__2166 (
            .O(N__21025),
            .I(N__21022));
    LocalMux I__2165 (
            .O(N__21022),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__2164 (
            .O(N__21019),
            .I(N__21016));
    LocalMux I__2163 (
            .O(N__21016),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__2162 (
            .O(N__21013),
            .I(N__21008));
    InMux I__2161 (
            .O(N__21012),
            .I(N__21005));
    InMux I__2160 (
            .O(N__21011),
            .I(N__21002));
    LocalMux I__2159 (
            .O(N__21008),
            .I(N__20997));
    LocalMux I__2158 (
            .O(N__21005),
            .I(N__20997));
    LocalMux I__2157 (
            .O(N__21002),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__2156 (
            .O(N__20997),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__2155 (
            .O(N__20992),
            .I(N__20989));
    LocalMux I__2154 (
            .O(N__20989),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__2153 (
            .O(N__20986),
            .I(N__20981));
    InMux I__2152 (
            .O(N__20985),
            .I(N__20978));
    InMux I__2151 (
            .O(N__20984),
            .I(N__20975));
    LocalMux I__2150 (
            .O(N__20981),
            .I(N__20972));
    LocalMux I__2149 (
            .O(N__20978),
            .I(N__20969));
    LocalMux I__2148 (
            .O(N__20975),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2147 (
            .O(N__20972),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2146 (
            .O(N__20969),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    CascadeMux I__2145 (
            .O(N__20962),
            .I(N__20959));
    InMux I__2144 (
            .O(N__20959),
            .I(N__20956));
    LocalMux I__2143 (
            .O(N__20956),
            .I(\pwm_generator_inst.counter_i_7 ));
    InMux I__2142 (
            .O(N__20953),
            .I(N__20949));
    InMux I__2141 (
            .O(N__20952),
            .I(N__20945));
    LocalMux I__2140 (
            .O(N__20949),
            .I(N__20942));
    InMux I__2139 (
            .O(N__20948),
            .I(N__20939));
    LocalMux I__2138 (
            .O(N__20945),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__2137 (
            .O(N__20942),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2136 (
            .O(N__20939),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2135 (
            .O(N__20932),
            .I(N__20929));
    LocalMux I__2134 (
            .O(N__20929),
            .I(\pwm_generator_inst.counter_i_8 ));
    InMux I__2133 (
            .O(N__20926),
            .I(N__20922));
    InMux I__2132 (
            .O(N__20925),
            .I(N__20918));
    LocalMux I__2131 (
            .O(N__20922),
            .I(N__20915));
    InMux I__2130 (
            .O(N__20921),
            .I(N__20912));
    LocalMux I__2129 (
            .O(N__20918),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__2128 (
            .O(N__20915),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2127 (
            .O(N__20912),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__2126 (
            .O(N__20905),
            .I(N__20902));
    LocalMux I__2125 (
            .O(N__20902),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2124 (
            .O(N__20899),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2123 (
            .O(N__20896),
            .I(N__20893));
    LocalMux I__2122 (
            .O(N__20893),
            .I(N__20890));
    Span4Mux_s3_v I__2121 (
            .O(N__20890),
            .I(N__20887));
    Span4Mux_v I__2120 (
            .O(N__20887),
            .I(N__20884));
    Sp12to4 I__2119 (
            .O(N__20884),
            .I(N__20881));
    Span12Mux_h I__2118 (
            .O(N__20881),
            .I(N__20878));
    Odrv12 I__2117 (
            .O(N__20878),
            .I(pwm_output_c));
    InMux I__2116 (
            .O(N__20875),
            .I(N__20872));
    LocalMux I__2115 (
            .O(N__20872),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    InMux I__2114 (
            .O(N__20869),
            .I(N__20866));
    LocalMux I__2113 (
            .O(N__20866),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__2112 (
            .O(N__20863),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    InMux I__2111 (
            .O(N__20860),
            .I(N__20857));
    LocalMux I__2110 (
            .O(N__20857),
            .I(N__20854));
    Odrv4 I__2109 (
            .O(N__20854),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    InMux I__2108 (
            .O(N__20851),
            .I(N__20848));
    LocalMux I__2107 (
            .O(N__20848),
            .I(N__20845));
    Odrv4 I__2106 (
            .O(N__20845),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1 ));
    InMux I__2105 (
            .O(N__20842),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__2104 (
            .O(N__20839),
            .I(N__20835));
    InMux I__2103 (
            .O(N__20838),
            .I(N__20831));
    LocalMux I__2102 (
            .O(N__20835),
            .I(N__20828));
    InMux I__2101 (
            .O(N__20834),
            .I(N__20825));
    LocalMux I__2100 (
            .O(N__20831),
            .I(N__20820));
    Span4Mux_h I__2099 (
            .O(N__20828),
            .I(N__20820));
    LocalMux I__2098 (
            .O(N__20825),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__2097 (
            .O(N__20820),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2096 (
            .O(N__20815),
            .I(N__20812));
    LocalMux I__2095 (
            .O(N__20812),
            .I(\pwm_generator_inst.counter_i_0 ));
    InMux I__2094 (
            .O(N__20809),
            .I(N__20804));
    InMux I__2093 (
            .O(N__20808),
            .I(N__20801));
    InMux I__2092 (
            .O(N__20807),
            .I(N__20798));
    LocalMux I__2091 (
            .O(N__20804),
            .I(N__20793));
    LocalMux I__2090 (
            .O(N__20801),
            .I(N__20793));
    LocalMux I__2089 (
            .O(N__20798),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__2088 (
            .O(N__20793),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__2087 (
            .O(N__20788),
            .I(N__20785));
    LocalMux I__2086 (
            .O(N__20785),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__2085 (
            .O(N__20782),
            .I(N__20779));
    InMux I__2084 (
            .O(N__20779),
            .I(N__20776));
    LocalMux I__2083 (
            .O(N__20776),
            .I(N__20773));
    Odrv4 I__2082 (
            .O(N__20773),
            .I(\pwm_generator_inst.threshold_2 ));
    InMux I__2081 (
            .O(N__20770),
            .I(N__20766));
    InMux I__2080 (
            .O(N__20769),
            .I(N__20763));
    LocalMux I__2079 (
            .O(N__20766),
            .I(N__20757));
    LocalMux I__2078 (
            .O(N__20763),
            .I(N__20757));
    InMux I__2077 (
            .O(N__20762),
            .I(N__20754));
    Span4Mux_v I__2076 (
            .O(N__20757),
            .I(N__20751));
    LocalMux I__2075 (
            .O(N__20754),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__2074 (
            .O(N__20751),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2073 (
            .O(N__20746),
            .I(N__20743));
    LocalMux I__2072 (
            .O(N__20743),
            .I(\pwm_generator_inst.counter_i_2 ));
    InMux I__2071 (
            .O(N__20740),
            .I(N__20735));
    InMux I__2070 (
            .O(N__20739),
            .I(N__20732));
    InMux I__2069 (
            .O(N__20738),
            .I(N__20729));
    LocalMux I__2068 (
            .O(N__20735),
            .I(N__20724));
    LocalMux I__2067 (
            .O(N__20732),
            .I(N__20724));
    LocalMux I__2066 (
            .O(N__20729),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__2065 (
            .O(N__20724),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    CascadeMux I__2064 (
            .O(N__20719),
            .I(N__20716));
    InMux I__2063 (
            .O(N__20716),
            .I(N__20713));
    LocalMux I__2062 (
            .O(N__20713),
            .I(N__20710));
    Odrv4 I__2061 (
            .O(N__20710),
            .I(\pwm_generator_inst.threshold_3 ));
    InMux I__2060 (
            .O(N__20707),
            .I(N__20704));
    LocalMux I__2059 (
            .O(N__20704),
            .I(\pwm_generator_inst.counter_i_3 ));
    InMux I__2058 (
            .O(N__20701),
            .I(N__20696));
    InMux I__2057 (
            .O(N__20700),
            .I(N__20693));
    InMux I__2056 (
            .O(N__20699),
            .I(N__20690));
    LocalMux I__2055 (
            .O(N__20696),
            .I(N__20685));
    LocalMux I__2054 (
            .O(N__20693),
            .I(N__20685));
    LocalMux I__2053 (
            .O(N__20690),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__2052 (
            .O(N__20685),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__2051 (
            .O(N__20680),
            .I(N__20677));
    LocalMux I__2050 (
            .O(N__20677),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__2049 (
            .O(N__20674),
            .I(N__20669));
    InMux I__2048 (
            .O(N__20673),
            .I(N__20666));
    InMux I__2047 (
            .O(N__20672),
            .I(N__20663));
    LocalMux I__2046 (
            .O(N__20669),
            .I(N__20658));
    LocalMux I__2045 (
            .O(N__20666),
            .I(N__20658));
    LocalMux I__2044 (
            .O(N__20663),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__2043 (
            .O(N__20658),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2042 (
            .O(N__20653),
            .I(N__20650));
    LocalMux I__2041 (
            .O(N__20650),
            .I(\pwm_generator_inst.counter_i_5 ));
    InMux I__2040 (
            .O(N__20647),
            .I(N__20644));
    LocalMux I__2039 (
            .O(N__20644),
            .I(N__20641));
    Odrv4 I__2038 (
            .O(N__20641),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ));
    InMux I__2037 (
            .O(N__20638),
            .I(N__20635));
    LocalMux I__2036 (
            .O(N__20635),
            .I(N__20632));
    Odrv4 I__2035 (
            .O(N__20632),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ));
    InMux I__2034 (
            .O(N__20629),
            .I(N__20626));
    LocalMux I__2033 (
            .O(N__20626),
            .I(N__20623));
    Odrv4 I__2032 (
            .O(N__20623),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ));
    InMux I__2031 (
            .O(N__20620),
            .I(N__20617));
    LocalMux I__2030 (
            .O(N__20617),
            .I(N__20614));
    Odrv4 I__2029 (
            .O(N__20614),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0 ));
    InMux I__2028 (
            .O(N__20611),
            .I(N__20608));
    LocalMux I__2027 (
            .O(N__20608),
            .I(N__20605));
    Odrv4 I__2026 (
            .O(N__20605),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0 ));
    InMux I__2025 (
            .O(N__20602),
            .I(N__20599));
    LocalMux I__2024 (
            .O(N__20599),
            .I(N__20596));
    Odrv4 I__2023 (
            .O(N__20596),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0 ));
    InMux I__2022 (
            .O(N__20593),
            .I(N__20590));
    LocalMux I__2021 (
            .O(N__20590),
            .I(N__20587));
    Odrv4 I__2020 (
            .O(N__20587),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0 ));
    InMux I__2019 (
            .O(N__20584),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__2018 (
            .O(N__20581),
            .I(N__20578));
    LocalMux I__2017 (
            .O(N__20578),
            .I(N__20575));
    Span4Mux_s2_h I__2016 (
            .O(N__20575),
            .I(N__20572));
    Odrv4 I__2015 (
            .O(N__20572),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    CascadeMux I__2014 (
            .O(N__20569),
            .I(N__20566));
    InMux I__2013 (
            .O(N__20566),
            .I(N__20563));
    LocalMux I__2012 (
            .O(N__20563),
            .I(N__20560));
    Odrv4 I__2011 (
            .O(N__20560),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ));
    InMux I__2010 (
            .O(N__20557),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__2009 (
            .O(N__20554),
            .I(N__20551));
    LocalMux I__2008 (
            .O(N__20551),
            .I(N__20548));
    Odrv4 I__2007 (
            .O(N__20548),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ));
    InMux I__2006 (
            .O(N__20545),
            .I(N__20541));
    InMux I__2005 (
            .O(N__20544),
            .I(N__20538));
    LocalMux I__2004 (
            .O(N__20541),
            .I(N__20535));
    LocalMux I__2003 (
            .O(N__20538),
            .I(N__20532));
    Odrv12 I__2002 (
            .O(N__20535),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8 ));
    Odrv4 I__2001 (
            .O(N__20532),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8 ));
    InMux I__2000 (
            .O(N__20527),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    CascadeMux I__1999 (
            .O(N__20524),
            .I(N__20521));
    InMux I__1998 (
            .O(N__20521),
            .I(N__20518));
    LocalMux I__1997 (
            .O(N__20518),
            .I(N__20515));
    Odrv4 I__1996 (
            .O(N__20515),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ));
    InMux I__1995 (
            .O(N__20512),
            .I(N__20509));
    LocalMux I__1994 (
            .O(N__20509),
            .I(N__20505));
    InMux I__1993 (
            .O(N__20508),
            .I(N__20502));
    Odrv4 I__1992 (
            .O(N__20505),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8 ));
    LocalMux I__1991 (
            .O(N__20502),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8 ));
    InMux I__1990 (
            .O(N__20497),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__1989 (
            .O(N__20494),
            .I(N__20491));
    LocalMux I__1988 (
            .O(N__20491),
            .I(N__20488));
    Odrv4 I__1987 (
            .O(N__20488),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ));
    InMux I__1986 (
            .O(N__20485),
            .I(bfn_2_14_0_));
    InMux I__1985 (
            .O(N__20482),
            .I(N__20479));
    LocalMux I__1984 (
            .O(N__20479),
            .I(N__20476));
    Odrv4 I__1983 (
            .O(N__20476),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ));
    InMux I__1982 (
            .O(N__20473),
            .I(N__20470));
    LocalMux I__1981 (
            .O(N__20470),
            .I(N__20467));
    Odrv4 I__1980 (
            .O(N__20467),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ));
    InMux I__1979 (
            .O(N__20464),
            .I(N__20461));
    LocalMux I__1978 (
            .O(N__20461),
            .I(N__20458));
    Odrv4 I__1977 (
            .O(N__20458),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ));
    InMux I__1976 (
            .O(N__20455),
            .I(N__20452));
    LocalMux I__1975 (
            .O(N__20452),
            .I(N__20449));
    Odrv4 I__1974 (
            .O(N__20449),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ));
    InMux I__1973 (
            .O(N__20446),
            .I(N__20442));
    InMux I__1972 (
            .O(N__20445),
            .I(N__20439));
    LocalMux I__1971 (
            .O(N__20442),
            .I(N__20436));
    LocalMux I__1970 (
            .O(N__20439),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv4 I__1969 (
            .O(N__20436),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__1968 (
            .O(N__20431),
            .I(N__20428));
    LocalMux I__1967 (
            .O(N__20428),
            .I(N__20425));
    Odrv4 I__1966 (
            .O(N__20425),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    CascadeMux I__1965 (
            .O(N__20422),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12_cascade_ ));
    CascadeMux I__1964 (
            .O(N__20419),
            .I(N__20416));
    InMux I__1963 (
            .O(N__20416),
            .I(N__20412));
    InMux I__1962 (
            .O(N__20415),
            .I(N__20409));
    LocalMux I__1961 (
            .O(N__20412),
            .I(N__20406));
    LocalMux I__1960 (
            .O(N__20409),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    Odrv4 I__1959 (
            .O(N__20406),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    InMux I__1958 (
            .O(N__20401),
            .I(N__20398));
    LocalMux I__1957 (
            .O(N__20398),
            .I(N__20395));
    Odrv4 I__1956 (
            .O(N__20395),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    CascadeMux I__1955 (
            .O(N__20392),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13_cascade_ ));
    InMux I__1954 (
            .O(N__20389),
            .I(N__20385));
    InMux I__1953 (
            .O(N__20388),
            .I(N__20382));
    LocalMux I__1952 (
            .O(N__20385),
            .I(N__20379));
    LocalMux I__1951 (
            .O(N__20382),
            .I(N__20376));
    Span4Mux_v I__1950 (
            .O(N__20379),
            .I(N__20371));
    Span4Mux_v I__1949 (
            .O(N__20376),
            .I(N__20371));
    Odrv4 I__1948 (
            .O(N__20371),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__1947 (
            .O(N__20368),
            .I(N__20365));
    LocalMux I__1946 (
            .O(N__20365),
            .I(N__20362));
    Span4Mux_h I__1945 (
            .O(N__20362),
            .I(N__20359));
    Odrv4 I__1944 (
            .O(N__20359),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1943 (
            .O(N__20356),
            .I(N__20350));
    InMux I__1942 (
            .O(N__20355),
            .I(N__20350));
    LocalMux I__1941 (
            .O(N__20350),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__1940 (
            .O(N__20347),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__1939 (
            .O(N__20344),
            .I(N__20341));
    LocalMux I__1938 (
            .O(N__20341),
            .I(N__20338));
    Span4Mux_h I__1937 (
            .O(N__20338),
            .I(N__20335));
    Odrv4 I__1936 (
            .O(N__20335),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1935 (
            .O(N__20332),
            .I(N__20326));
    InMux I__1934 (
            .O(N__20331),
            .I(N__20326));
    LocalMux I__1933 (
            .O(N__20326),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    InMux I__1932 (
            .O(N__20323),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__1931 (
            .O(N__20320),
            .I(N__20317));
    LocalMux I__1930 (
            .O(N__20317),
            .I(N__20314));
    Span4Mux_h I__1929 (
            .O(N__20314),
            .I(N__20311));
    Odrv4 I__1928 (
            .O(N__20311),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1927 (
            .O(N__20308),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__1926 (
            .O(N__20305),
            .I(N__20302));
    LocalMux I__1925 (
            .O(N__20302),
            .I(N__20299));
    Odrv4 I__1924 (
            .O(N__20299),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__1923 (
            .O(N__20296),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    InMux I__1922 (
            .O(N__20293),
            .I(N__20289));
    InMux I__1921 (
            .O(N__20292),
            .I(N__20286));
    LocalMux I__1920 (
            .O(N__20289),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    LocalMux I__1919 (
            .O(N__20286),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    InMux I__1918 (
            .O(N__20281),
            .I(N__20275));
    InMux I__1917 (
            .O(N__20280),
            .I(N__20275));
    LocalMux I__1916 (
            .O(N__20275),
            .I(N__20272));
    Span4Mux_h I__1915 (
            .O(N__20272),
            .I(N__20269));
    Odrv4 I__1914 (
            .O(N__20269),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1913 (
            .O(N__20266),
            .I(N__20263));
    LocalMux I__1912 (
            .O(N__20263),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    CascadeMux I__1911 (
            .O(N__20260),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10_cascade_ ));
    InMux I__1910 (
            .O(N__20257),
            .I(N__20253));
    InMux I__1909 (
            .O(N__20256),
            .I(N__20250));
    LocalMux I__1908 (
            .O(N__20253),
            .I(N__20247));
    LocalMux I__1907 (
            .O(N__20250),
            .I(pwm_duty_input_1));
    Odrv4 I__1906 (
            .O(N__20247),
            .I(pwm_duty_input_1));
    InMux I__1905 (
            .O(N__20242),
            .I(N__20239));
    LocalMux I__1904 (
            .O(N__20239),
            .I(N__20235));
    InMux I__1903 (
            .O(N__20238),
            .I(N__20232));
    Span4Mux_s1_h I__1902 (
            .O(N__20235),
            .I(N__20229));
    LocalMux I__1901 (
            .O(N__20232),
            .I(pwm_duty_input_0));
    Odrv4 I__1900 (
            .O(N__20229),
            .I(pwm_duty_input_0));
    InMux I__1899 (
            .O(N__20224),
            .I(N__20221));
    LocalMux I__1898 (
            .O(N__20221),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__1897 (
            .O(N__20218),
            .I(N__20213));
    InMux I__1896 (
            .O(N__20217),
            .I(N__20208));
    InMux I__1895 (
            .O(N__20216),
            .I(N__20208));
    LocalMux I__1894 (
            .O(N__20213),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    LocalMux I__1893 (
            .O(N__20208),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__1892 (
            .O(N__20203),
            .I(N__20200));
    LocalMux I__1891 (
            .O(N__20200),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__1890 (
            .O(N__20197),
            .I(N__20193));
    InMux I__1889 (
            .O(N__20196),
            .I(N__20189));
    LocalMux I__1888 (
            .O(N__20193),
            .I(N__20186));
    InMux I__1887 (
            .O(N__20192),
            .I(N__20183));
    LocalMux I__1886 (
            .O(N__20189),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    Odrv4 I__1885 (
            .O(N__20186),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__1884 (
            .O(N__20183),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    InMux I__1883 (
            .O(N__20176),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    InMux I__1882 (
            .O(N__20173),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__1881 (
            .O(N__20170),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__1880 (
            .O(N__20167),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    InMux I__1879 (
            .O(N__20164),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    InMux I__1878 (
            .O(N__20161),
            .I(bfn_2_10_0_));
    InMux I__1877 (
            .O(N__20158),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__1876 (
            .O(N__20155),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__1875 (
            .O(N__20152),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__1874 (
            .O(N__20149),
            .I(N__20146));
    LocalMux I__1873 (
            .O(N__20146),
            .I(N__20143));
    Span4Mux_v I__1872 (
            .O(N__20143),
            .I(N__20140));
    Odrv4 I__1871 (
            .O(N__20140),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1870 (
            .O(N__20137),
            .I(N__20134));
    LocalMux I__1869 (
            .O(N__20134),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__1868 (
            .O(N__20131),
            .I(N__20128));
    LocalMux I__1867 (
            .O(N__20128),
            .I(N__20125));
    Span4Mux_h I__1866 (
            .O(N__20125),
            .I(N__20122));
    Odrv4 I__1865 (
            .O(N__20122),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1864 (
            .O(N__20119),
            .I(N__20116));
    LocalMux I__1863 (
            .O(N__20116),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    InMux I__1862 (
            .O(N__20113),
            .I(N__20110));
    LocalMux I__1861 (
            .O(N__20110),
            .I(N__20107));
    Span4Mux_h I__1860 (
            .O(N__20107),
            .I(N__20104));
    Odrv4 I__1859 (
            .O(N__20104),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1858 (
            .O(N__20101),
            .I(N__20098));
    LocalMux I__1857 (
            .O(N__20098),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__1856 (
            .O(N__20095),
            .I(N__20092));
    LocalMux I__1855 (
            .O(N__20092),
            .I(N__20089));
    Span4Mux_h I__1854 (
            .O(N__20089),
            .I(N__20086));
    Odrv4 I__1853 (
            .O(N__20086),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1852 (
            .O(N__20083),
            .I(N__20080));
    LocalMux I__1851 (
            .O(N__20080),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__1850 (
            .O(N__20077),
            .I(N__20074));
    LocalMux I__1849 (
            .O(N__20074),
            .I(N__20071));
    Span4Mux_h I__1848 (
            .O(N__20071),
            .I(N__20068));
    Odrv4 I__1847 (
            .O(N__20068),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1846 (
            .O(N__20065),
            .I(N__20062));
    LocalMux I__1845 (
            .O(N__20062),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__1844 (
            .O(N__20059),
            .I(N__20056));
    LocalMux I__1843 (
            .O(N__20056),
            .I(N__20053));
    Span4Mux_h I__1842 (
            .O(N__20053),
            .I(N__20050));
    Odrv4 I__1841 (
            .O(N__20050),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1840 (
            .O(N__20047),
            .I(N__20044));
    LocalMux I__1839 (
            .O(N__20044),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__1838 (
            .O(N__20041),
            .I(N__20038));
    LocalMux I__1837 (
            .O(N__20038),
            .I(N__20035));
    Span4Mux_h I__1836 (
            .O(N__20035),
            .I(N__20032));
    Odrv4 I__1835 (
            .O(N__20032),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1834 (
            .O(N__20029),
            .I(N__20026));
    LocalMux I__1833 (
            .O(N__20026),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__1832 (
            .O(N__20023),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    InMux I__1831 (
            .O(N__20020),
            .I(bfn_2_6_0_));
    InMux I__1830 (
            .O(N__20017),
            .I(\pwm_generator_inst.counter_cry_8 ));
    CascadeMux I__1829 (
            .O(N__20014),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    CascadeMux I__1828 (
            .O(N__20011),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__1827 (
            .O(N__20008),
            .I(N__19990));
    InMux I__1826 (
            .O(N__20007),
            .I(N__19990));
    InMux I__1825 (
            .O(N__20006),
            .I(N__19990));
    InMux I__1824 (
            .O(N__20005),
            .I(N__19990));
    InMux I__1823 (
            .O(N__20004),
            .I(N__19981));
    InMux I__1822 (
            .O(N__20003),
            .I(N__19981));
    InMux I__1821 (
            .O(N__20002),
            .I(N__19981));
    InMux I__1820 (
            .O(N__20001),
            .I(N__19981));
    InMux I__1819 (
            .O(N__20000),
            .I(N__19976));
    InMux I__1818 (
            .O(N__19999),
            .I(N__19976));
    LocalMux I__1817 (
            .O(N__19990),
            .I(N__19971));
    LocalMux I__1816 (
            .O(N__19981),
            .I(N__19971));
    LocalMux I__1815 (
            .O(N__19976),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__1814 (
            .O(N__19971),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__1813 (
            .O(N__19966),
            .I(N__19963));
    LocalMux I__1812 (
            .O(N__19963),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    InMux I__1811 (
            .O(N__19960),
            .I(N__19957));
    LocalMux I__1810 (
            .O(N__19957),
            .I(N__19954));
    Span4Mux_h I__1809 (
            .O(N__19954),
            .I(N__19951));
    Odrv4 I__1808 (
            .O(N__19951),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1807 (
            .O(N__19948),
            .I(N__19945));
    LocalMux I__1806 (
            .O(N__19945),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__1805 (
            .O(N__19942),
            .I(N__19939));
    LocalMux I__1804 (
            .O(N__19939),
            .I(N__19936));
    Span4Mux_h I__1803 (
            .O(N__19936),
            .I(N__19933));
    Odrv4 I__1802 (
            .O(N__19933),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1801 (
            .O(N__19930),
            .I(N__19927));
    LocalMux I__1800 (
            .O(N__19927),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__1799 (
            .O(N__19924),
            .I(N__19921));
    LocalMux I__1798 (
            .O(N__19921),
            .I(N__19918));
    Span4Mux_v I__1797 (
            .O(N__19918),
            .I(N__19915));
    Odrv4 I__1796 (
            .O(N__19915),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1795 (
            .O(N__19912),
            .I(N__19909));
    LocalMux I__1794 (
            .O(N__19909),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__1793 (
            .O(N__19906),
            .I(N__19903));
    LocalMux I__1792 (
            .O(N__19903),
            .I(un7_start_stop_0_a2));
    InMux I__1791 (
            .O(N__19900),
            .I(bfn_2_5_0_));
    InMux I__1790 (
            .O(N__19897),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__1789 (
            .O(N__19894),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__1788 (
            .O(N__19891),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__1787 (
            .O(N__19888),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__1786 (
            .O(N__19885),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__1785 (
            .O(N__19882),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__1784 (
            .O(N__19879),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__1783 (
            .O(N__19876),
            .I(N__19873));
    LocalMux I__1782 (
            .O(N__19873),
            .I(N__19870));
    Span4Mux_v I__1781 (
            .O(N__19870),
            .I(N__19867));
    Odrv4 I__1780 (
            .O(N__19867),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__1779 (
            .O(N__19864),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    InMux I__1778 (
            .O(N__19861),
            .I(N__19858));
    LocalMux I__1777 (
            .O(N__19858),
            .I(N__19855));
    Span4Mux_v I__1776 (
            .O(N__19855),
            .I(N__19852));
    Odrv4 I__1775 (
            .O(N__19852),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__1774 (
            .O(N__19849),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    InMux I__1773 (
            .O(N__19846),
            .I(N__19843));
    LocalMux I__1772 (
            .O(N__19843),
            .I(N__19840));
    Span4Mux_v I__1771 (
            .O(N__19840),
            .I(N__19837));
    Odrv4 I__1770 (
            .O(N__19837),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    InMux I__1769 (
            .O(N__19834),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    InMux I__1768 (
            .O(N__19831),
            .I(N__19828));
    LocalMux I__1767 (
            .O(N__19828),
            .I(N__19825));
    Span4Mux_v I__1766 (
            .O(N__19825),
            .I(N__19822));
    Odrv4 I__1765 (
            .O(N__19822),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__1764 (
            .O(N__19819),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    CascadeMux I__1763 (
            .O(N__19816),
            .I(N__19813));
    InMux I__1762 (
            .O(N__19813),
            .I(N__19810));
    LocalMux I__1761 (
            .O(N__19810),
            .I(N__19807));
    Span12Mux_v I__1760 (
            .O(N__19807),
            .I(N__19804));
    Odrv12 I__1759 (
            .O(N__19804),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    InMux I__1758 (
            .O(N__19801),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__1757 (
            .O(N__19798),
            .I(bfn_1_13_0_));
    InMux I__1756 (
            .O(N__19795),
            .I(N__19792));
    LocalMux I__1755 (
            .O(N__19792),
            .I(N__19789));
    Span4Mux_v I__1754 (
            .O(N__19789),
            .I(N__19786));
    Odrv4 I__1753 (
            .O(N__19786),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__1752 (
            .O(N__19783),
            .I(N__19780));
    LocalMux I__1751 (
            .O(N__19780),
            .I(N__19777));
    Span4Mux_v I__1750 (
            .O(N__19777),
            .I(N__19769));
    CascadeMux I__1749 (
            .O(N__19776),
            .I(N__19765));
    CascadeMux I__1748 (
            .O(N__19775),
            .I(N__19762));
    CascadeMux I__1747 (
            .O(N__19774),
            .I(N__19758));
    CascadeMux I__1746 (
            .O(N__19773),
            .I(N__19755));
    CascadeMux I__1745 (
            .O(N__19772),
            .I(N__19752));
    Span4Mux_v I__1744 (
            .O(N__19769),
            .I(N__19749));
    InMux I__1743 (
            .O(N__19768),
            .I(N__19746));
    InMux I__1742 (
            .O(N__19765),
            .I(N__19741));
    InMux I__1741 (
            .O(N__19762),
            .I(N__19741));
    InMux I__1740 (
            .O(N__19761),
            .I(N__19732));
    InMux I__1739 (
            .O(N__19758),
            .I(N__19732));
    InMux I__1738 (
            .O(N__19755),
            .I(N__19732));
    InMux I__1737 (
            .O(N__19752),
            .I(N__19732));
    Odrv4 I__1736 (
            .O(N__19749),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    LocalMux I__1735 (
            .O(N__19746),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    LocalMux I__1734 (
            .O(N__19741),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    LocalMux I__1733 (
            .O(N__19732),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    CascadeMux I__1732 (
            .O(N__19723),
            .I(N__19720));
    InMux I__1731 (
            .O(N__19720),
            .I(N__19717));
    LocalMux I__1730 (
            .O(N__19717),
            .I(N__19713));
    InMux I__1729 (
            .O(N__19716),
            .I(N__19710));
    Span4Mux_v I__1728 (
            .O(N__19713),
            .I(N__19707));
    LocalMux I__1727 (
            .O(N__19710),
            .I(N__19704));
    Odrv4 I__1726 (
            .O(N__19707),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    Odrv4 I__1725 (
            .O(N__19704),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    InMux I__1724 (
            .O(N__19699),
            .I(N__19696));
    LocalMux I__1723 (
            .O(N__19696),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__1722 (
            .O(N__19693),
            .I(N__19690));
    LocalMux I__1721 (
            .O(N__19690),
            .I(N_42_i_i));
    InMux I__1720 (
            .O(N__19687),
            .I(N__19684));
    LocalMux I__1719 (
            .O(N__19684),
            .I(N__19681));
    Span4Mux_v I__1718 (
            .O(N__19681),
            .I(N__19678));
    Odrv4 I__1717 (
            .O(N__19678),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__1716 (
            .O(N__19675),
            .I(N__19672));
    InMux I__1715 (
            .O(N__19672),
            .I(N__19669));
    LocalMux I__1714 (
            .O(N__19669),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    InMux I__1713 (
            .O(N__19666),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__1712 (
            .O(N__19663),
            .I(N__19660));
    LocalMux I__1711 (
            .O(N__19660),
            .I(N__19657));
    Span4Mux_v I__1710 (
            .O(N__19657),
            .I(N__19654));
    Odrv4 I__1709 (
            .O(N__19654),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    CascadeMux I__1708 (
            .O(N__19651),
            .I(N__19648));
    InMux I__1707 (
            .O(N__19648),
            .I(N__19645));
    LocalMux I__1706 (
            .O(N__19645),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__1705 (
            .O(N__19642),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__1704 (
            .O(N__19639),
            .I(N__19636));
    LocalMux I__1703 (
            .O(N__19636),
            .I(N__19633));
    Span4Mux_v I__1702 (
            .O(N__19633),
            .I(N__19630));
    Odrv4 I__1701 (
            .O(N__19630),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__1700 (
            .O(N__19627),
            .I(N__19624));
    InMux I__1699 (
            .O(N__19624),
            .I(N__19621));
    LocalMux I__1698 (
            .O(N__19621),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    InMux I__1697 (
            .O(N__19618),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__1696 (
            .O(N__19615),
            .I(N__19612));
    LocalMux I__1695 (
            .O(N__19612),
            .I(N__19609));
    Span4Mux_v I__1694 (
            .O(N__19609),
            .I(N__19606));
    Odrv4 I__1693 (
            .O(N__19606),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    CascadeMux I__1692 (
            .O(N__19603),
            .I(N__19600));
    InMux I__1691 (
            .O(N__19600),
            .I(N__19597));
    LocalMux I__1690 (
            .O(N__19597),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    InMux I__1689 (
            .O(N__19594),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__1688 (
            .O(N__19591),
            .I(N__19588));
    LocalMux I__1687 (
            .O(N__19588),
            .I(N__19585));
    Span4Mux_v I__1686 (
            .O(N__19585),
            .I(N__19582));
    Odrv4 I__1685 (
            .O(N__19582),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    CascadeMux I__1684 (
            .O(N__19579),
            .I(N__19576));
    InMux I__1683 (
            .O(N__19576),
            .I(N__19573));
    LocalMux I__1682 (
            .O(N__19573),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    InMux I__1681 (
            .O(N__19570),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__1680 (
            .O(N__19567),
            .I(N__19564));
    LocalMux I__1679 (
            .O(N__19564),
            .I(N__19561));
    Span4Mux_v I__1678 (
            .O(N__19561),
            .I(N__19558));
    Odrv4 I__1677 (
            .O(N__19558),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    CascadeMux I__1676 (
            .O(N__19555),
            .I(N__19552));
    InMux I__1675 (
            .O(N__19552),
            .I(N__19549));
    LocalMux I__1674 (
            .O(N__19549),
            .I(N__19546));
    Odrv4 I__1673 (
            .O(N__19546),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    InMux I__1672 (
            .O(N__19543),
            .I(bfn_1_12_0_));
    InMux I__1671 (
            .O(N__19540),
            .I(N__19537));
    LocalMux I__1670 (
            .O(N__19537),
            .I(N__19534));
    Span4Mux_v I__1669 (
            .O(N__19534),
            .I(N__19531));
    Odrv4 I__1668 (
            .O(N__19531),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    CascadeMux I__1667 (
            .O(N__19528),
            .I(N__19525));
    InMux I__1666 (
            .O(N__19525),
            .I(N__19522));
    LocalMux I__1665 (
            .O(N__19522),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    InMux I__1664 (
            .O(N__19519),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    InMux I__1663 (
            .O(N__19516),
            .I(N__19513));
    LocalMux I__1662 (
            .O(N__19513),
            .I(N__19510));
    Span4Mux_v I__1661 (
            .O(N__19510),
            .I(N__19507));
    Odrv4 I__1660 (
            .O(N__19507),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__1659 (
            .O(N__19504),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    InMux I__1658 (
            .O(N__19501),
            .I(N__19498));
    LocalMux I__1657 (
            .O(N__19498),
            .I(N__19495));
    Span4Mux_v I__1656 (
            .O(N__19495),
            .I(N__19492));
    Odrv4 I__1655 (
            .O(N__19492),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__1654 (
            .O(N__19489),
            .I(N__19486));
    InMux I__1653 (
            .O(N__19486),
            .I(N__19483));
    LocalMux I__1652 (
            .O(N__19483),
            .I(N__19480));
    Odrv4 I__1651 (
            .O(N__19480),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__1650 (
            .O(N__19477),
            .I(N__19474));
    LocalMux I__1649 (
            .O(N__19474),
            .I(N__19471));
    Span4Mux_v I__1648 (
            .O(N__19471),
            .I(N__19468));
    Odrv4 I__1647 (
            .O(N__19468),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__1646 (
            .O(N__19465),
            .I(N__19462));
    InMux I__1645 (
            .O(N__19462),
            .I(N__19459));
    LocalMux I__1644 (
            .O(N__19459),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    InMux I__1643 (
            .O(N__19456),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__1642 (
            .O(N__19453),
            .I(N__19450));
    LocalMux I__1641 (
            .O(N__19450),
            .I(N__19447));
    Span4Mux_v I__1640 (
            .O(N__19447),
            .I(N__19444));
    Odrv4 I__1639 (
            .O(N__19444),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__1638 (
            .O(N__19441),
            .I(N__19438));
    InMux I__1637 (
            .O(N__19438),
            .I(N__19435));
    LocalMux I__1636 (
            .O(N__19435),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__1635 (
            .O(N__19432),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    IoInMux I__1634 (
            .O(N__19429),
            .I(N__19426));
    LocalMux I__1633 (
            .O(N__19426),
            .I(N__19423));
    Span4Mux_s3_v I__1632 (
            .O(N__19423),
            .I(N__19420));
    Span4Mux_h I__1631 (
            .O(N__19420),
            .I(N__19417));
    Sp12to4 I__1630 (
            .O(N__19417),
            .I(N__19414));
    Span12Mux_v I__1629 (
            .O(N__19414),
            .I(N__19411));
    Span12Mux_v I__1628 (
            .O(N__19411),
            .I(N__19408));
    Odrv12 I__1627 (
            .O(N__19408),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1626 (
            .O(N__19405),
            .I(N__19402));
    LocalMux I__1625 (
            .O(N__19402),
            .I(N__19399));
    IoSpan4Mux I__1624 (
            .O(N__19399),
            .I(N__19396));
    IoSpan4Mux I__1623 (
            .O(N__19396),
            .I(N__19393));
    Odrv4 I__1622 (
            .O(N__19393),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_10_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_25_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_10_25_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_3_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_10_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_3_10_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_3_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_7_0_));
    defparam IN_MUX_bfv_3_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_8_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_3_8_0_));
    defparam IN_MUX_bfv_2_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_5_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_13_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_14_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_13_14_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_11_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_21_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_11_21_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_17_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_17_8_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_15_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_22_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_15_22_0_));
    defparam IN_MUX_bfv_15_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_23_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_15_23_0_));
    defparam IN_MUX_bfv_15_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_24_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_15_24_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_7_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_7_21_0_));
    defparam IN_MUX_bfv_7_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_7_22_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_8_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_23_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_8_23_0_));
    defparam IN_MUX_bfv_8_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_24_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_8_24_0_));
    defparam IN_MUX_bfv_13_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_4_0_));
    defparam IN_MUX_bfv_13_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_5_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .carryinitout(bfn_13_5_0_));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_12_10_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19429),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19405),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__26158),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_hc_timer.N_397_i_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__34831),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_166_i_g ));
    ICE_GB \delay_measurement_inst.delay_tr_timer.running_RNICNBI_0  (
            .USERSIGNALTOGLOBALBUFFER(N__28960),
            .GLOBALBUFFEROUTPUT(\delay_measurement_inst.delay_tr_timer.N_399_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__28304),
            .CLKHFEN(N__28308),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__28315),
            .RGB2PWM(N__19693),
            .RGB1(rgb_g),
            .CURREN(N__28309),
            .RGB2(rgb_b),
            .RGB1PWM(N__19906),
            .RGB0PWM(N__49588),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_4_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_4_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_4_6  (
            .in0(N__19783),
            .in1(N__19716),
            .in2(_gnd_net_),
            .in3(N__21378),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23176),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49977),
            .ce(),
            .sr(N__49496));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_9_5 .LUT_INIT=16'b1111010001010100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_9_5  (
            .in0(N__23175),
            .in1(N__22123),
            .in2(N__22578),
            .in3(N__22358),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49975),
            .ce(),
            .sr(N__49516));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_0 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_10_0  (
            .in0(N__21768),
            .in1(N__22435),
            .in2(N__22182),
            .in3(N__22266),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(),
            .sr(N__49520));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_2 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_10_2  (
            .in0(N__22420),
            .in1(N__21769),
            .in2(N__22183),
            .in3(N__22267),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(),
            .sr(N__49520));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_10_3  (
            .in0(N__21253),
            .in1(N__22355),
            .in2(N__21235),
            .in3(N__22696),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(),
            .sr(N__49520));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_4 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_10_4  (
            .in0(N__23169),
            .in1(N__22615),
            .in2(N__22359),
            .in3(N__22121),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(),
            .sr(N__49520));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_5 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_10_5  (
            .in0(N__22119),
            .in1(N__23168),
            .in2(N__22657),
            .in3(N__22356),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(),
            .sr(N__49520));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_6 .LUT_INIT=16'b1101010111000100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_10_6  (
            .in0(N__23170),
            .in1(N__22543),
            .in2(N__22360),
            .in3(N__22122),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(),
            .sr(N__49520));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7 .LUT_INIT=16'b1111001000110010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_10_7  (
            .in0(N__22120),
            .in1(N__23171),
            .in2(N__22507),
            .in3(N__22357),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49973),
            .ce(),
            .sr(N__49520));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_1_11_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_1_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__19501),
            .in2(N__19489),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_11_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__19477),
            .in2(N__19465),
            .in3(N__19456),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_11_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__19453),
            .in2(N__19441),
            .in3(N__19432),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_11_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__19687),
            .in2(N__19675),
            .in3(N__19666),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_11_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__19663),
            .in2(N__19651),
            .in3(N__19642),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_11_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__19639),
            .in2(N__19627),
            .in3(N__19618),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_11_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__19615),
            .in2(N__19603),
            .in3(N__19594),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_11_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__19591),
            .in2(N__19579),
            .in3(N__19570),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__19567),
            .in2(N__19555),
            .in3(N__19543),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__19540),
            .in2(N__19528),
            .in3(N__19519),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__19516),
            .in2(N__19772),
            .in3(N__19504),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__19876),
            .in2(N__19775),
            .in3(N__19864),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_12_s_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__19861),
            .in2(N__19773),
            .in3(N__19849),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_12_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_13_s_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__19846),
            .in2(N__19776),
            .in3(N__19834),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_13_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_14_s_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__19831),
            .in2(N__19774),
            .in3(N__19819),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_14_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_s_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(N__19761),
            .in2(N__19816),
            .in3(N__19801),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_13_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHR5_LC_1_13_0  (
            .in0(N__20581),
            .in1(N__19699),
            .in2(_gnd_net_),
            .in3(N__19798),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNIFHRZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_5 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_13_5  (
            .in0(N__19795),
            .in1(N__19768),
            .in2(N__19723),
            .in3(N__21411),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.N_42_i_i_LC_1_29_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.N_42_i_i_LC_1_29_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.N_42_i_i_LC_1_29_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \phase_controller_inst1.N_42_i_i_LC_1_29_7  (
            .in0(N__33156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49586),
            .lcout(N_42_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_5  (
            .in0(N__33160),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49587),
            .lcout(un7_start_stop_0_a2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_2_5_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_2_5_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_2_5_0  (
            .in0(N__20005),
            .in1(N__20834),
            .in2(_gnd_net_),
            .in3(N__19900),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_5_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__49978),
            .ce(),
            .sr(N__49483));
    defparam \pwm_generator_inst.counter_1_LC_2_5_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_2_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_2_5_1  (
            .in0(N__20001),
            .in1(N__20807),
            .in2(_gnd_net_),
            .in3(N__19897),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__49978),
            .ce(),
            .sr(N__49483));
    defparam \pwm_generator_inst.counter_2_LC_2_5_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_2_5_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_2_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_2_5_2  (
            .in0(N__20006),
            .in1(N__20762),
            .in2(_gnd_net_),
            .in3(N__19894),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__49978),
            .ce(),
            .sr(N__49483));
    defparam \pwm_generator_inst.counter_3_LC_2_5_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_2_5_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_2_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_2_5_3  (
            .in0(N__20002),
            .in1(N__20738),
            .in2(_gnd_net_),
            .in3(N__19891),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__49978),
            .ce(),
            .sr(N__49483));
    defparam \pwm_generator_inst.counter_4_LC_2_5_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_2_5_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_2_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_2_5_4  (
            .in0(N__20007),
            .in1(N__20699),
            .in2(_gnd_net_),
            .in3(N__19888),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__49978),
            .ce(),
            .sr(N__49483));
    defparam \pwm_generator_inst.counter_5_LC_2_5_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_2_5_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_2_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_2_5_5  (
            .in0(N__20003),
            .in1(N__20672),
            .in2(_gnd_net_),
            .in3(N__19885),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__49978),
            .ce(),
            .sr(N__49483));
    defparam \pwm_generator_inst.counter_6_LC_2_5_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_2_5_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_2_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_2_5_6  (
            .in0(N__20008),
            .in1(N__21011),
            .in2(_gnd_net_),
            .in3(N__19882),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__49978),
            .ce(),
            .sr(N__49483));
    defparam \pwm_generator_inst.counter_7_LC_2_5_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_2_5_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_2_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_2_5_7  (
            .in0(N__20004),
            .in1(N__20984),
            .in2(_gnd_net_),
            .in3(N__19879),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__49978),
            .ce(),
            .sr(N__49483));
    defparam \pwm_generator_inst.counter_8_LC_2_6_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_2_6_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_2_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_2_6_0  (
            .in0(N__20000),
            .in1(N__20952),
            .in2(_gnd_net_),
            .in3(N__20020),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__49976),
            .ce(),
            .sr(N__49490));
    defparam \pwm_generator_inst.counter_9_LC_2_6_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_2_6_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_2_6_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_2_6_1  (
            .in0(N__20925),
            .in1(N__19999),
            .in2(_gnd_net_),
            .in3(N__20017),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49976),
            .ce(),
            .sr(N__49490));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_2_7_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_2_7_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__20838),
            .in2(_gnd_net_),
            .in3(N__20770),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_2_7_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_2_7_2 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_2_7_2  (
            .in0(N__20701),
            .in1(N__20740),
            .in2(N__20014),
            .in3(N__20809),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_2_7_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_2_7_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_2_7_3  (
            .in0(N__19966),
            .in1(N__21013),
            .in2(N__20011),
            .in3(N__20674),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_2_7_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_2_7_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_2_7_4  (
            .in0(N__20985),
            .in1(N__20921),
            .in2(_gnd_net_),
            .in3(N__20948),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__19948),
            .in2(_gnd_net_),
            .in3(N__19960),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__19930),
            .in2(_gnd_net_),
            .in3(N__19942),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_8_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__19912),
            .in2(_gnd_net_),
            .in3(N__19924),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_8_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_8_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_8_3  (
            .in0(N__20149),
            .in1(N__20137),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_8_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__20119),
            .in2(_gnd_net_),
            .in3(N__20131),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_8_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__20101),
            .in2(_gnd_net_),
            .in3(N__20113),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_8_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__20083),
            .in2(_gnd_net_),
            .in3(N__20095),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_8_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(N__20065),
            .in2(_gnd_net_),
            .in3(N__20077),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__20047),
            .in2(_gnd_net_),
            .in3(N__20059),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__20029),
            .in2(_gnd_net_),
            .in3(N__20041),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__20292),
            .in2(_gnd_net_),
            .in3(N__20023),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_2_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_2_9_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNI5VQP_LC_2_9_3  (
            .in0(N__21998),
            .in1(N__20389),
            .in2(_gnd_net_),
            .in3(N__20176),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__20446),
            .in2(_gnd_net_),
            .in3(N__20173),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20419),
            .in3(N__20170),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__21204),
            .in2(_gnd_net_),
            .in3(N__20167),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__22059),
            .in2(_gnd_net_),
            .in3(N__20164),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__21041),
            .in2(_gnd_net_),
            .in3(N__20161),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_10_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__20216),
            .in2(_gnd_net_),
            .in3(N__20158),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_10_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__20197),
            .in2(_gnd_net_),
            .in3(N__20155),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_10_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20152),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_10_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_2_10_4  (
            .in0(N__20293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20280),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_2_10_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_2_10_5 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIT6OT_LC_2_10_5  (
            .in0(N__20281),
            .in1(N__20266),
            .in2(N__20260),
            .in3(N__21981),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_10_6  (
            .in0(N__21744),
            .in1(N__20256),
            .in2(_gnd_net_),
            .in3(N__20238),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_2_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_2_10_7 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNI6DBN_LC_2_10_7  (
            .in0(N__20224),
            .in1(N__20217),
            .in2(N__22003),
            .in3(N__20545),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_11_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__20218),
            .in2(_gnd_net_),
            .in3(N__20544),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_2_11_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_2_11_4 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNI9JEN_LC_2_11_4  (
            .in0(N__20192),
            .in1(N__20512),
            .in2(N__22004),
            .in3(N__20203),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_11_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_11_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__21063),
            .in2(_gnd_net_),
            .in3(N__21045),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_12_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_12_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_12_0  (
            .in0(N__20508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20196),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_12_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_12_1  (
            .in0(N__22058),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22026),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_12_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_12_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__20355),
            .in2(_gnd_net_),
            .in3(N__20445),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_2_12_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_2_12_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNIBKRQ_LC_2_12_4  (
            .in0(N__20356),
            .in1(N__20431),
            .in2(N__20422),
            .in3(N__21967),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_2_12_5  (
            .in0(N__20415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20331),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_2_12_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_2_12_6 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIDOTQ_LC_2_12_6  (
            .in0(N__20332),
            .in1(N__20401),
            .in2(N__20392),
            .in3(N__21968),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__20388),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__20368),
            .in2(_gnd_net_),
            .in3(N__20347),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__20344),
            .in2(_gnd_net_),
            .in3(N__20323),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__20320),
            .in2(_gnd_net_),
            .in3(N__20308),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__20305),
            .in2(_gnd_net_),
            .in3(N__20296),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIM5E8_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__28277),
            .in2(N__20569),
            .in3(N__20557),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIM5EZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIO9G8_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__20554),
            .in2(N__28310),
            .in3(N__20527),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIO9GZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIQDI8_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__28281),
            .in2(N__20524),
            .in3(N__20497),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIQDIZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNISHK8_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__20494),
            .in2(_gnd_net_),
            .in3(N__20485),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNISHKZ0Z8 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__20482),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__20473),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__20464),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__20455),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__20647),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__20638),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__20629),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__20620),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__20611),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__20602),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__20593),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_15_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20584),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_3_6_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_3_6_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_3_6_5 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIS7985_LC_3_6_5  (
            .in0(N__21598),
            .in1(N__20851),
            .in2(N__21428),
            .in3(N__21813),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_6_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_6_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_6_7 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIVDC85_LC_3_6_7  (
            .in0(N__21599),
            .in1(N__21124),
            .in2(N__21429),
            .in3(N__21814),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_7_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_7_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_7_0  (
            .in0(_gnd_net_),
            .in1(N__20815),
            .in2(N__21145),
            .in3(N__20839),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_3_7_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_7_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_7_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_7_1  (
            .in0(_gnd_net_),
            .in1(N__20788),
            .in2(N__21472),
            .in3(N__20808),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_7_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_7_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_7_2  (
            .in0(_gnd_net_),
            .in1(N__20746),
            .in2(N__20782),
            .in3(N__20769),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_7_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_7_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_7_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_7_3  (
            .in0(N__20739),
            .in1(N__20707),
            .in2(N__20719),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_7_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_7_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_7_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_7_4  (
            .in0(N__20700),
            .in1(N__20680),
            .in2(N__21487),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_7_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_7_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_7_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_7_5  (
            .in0(N__20673),
            .in1(N__20653),
            .in2(N__21523),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_7_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_7_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_7_6  (
            .in0(N__21012),
            .in1(N__20992),
            .in2(N__21508),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_7_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_7_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_7_7  (
            .in0(_gnd_net_),
            .in1(N__21277),
            .in2(N__20962),
            .in3(N__20986),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_8_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_8_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_8_0  (
            .in0(N__20953),
            .in1(N__20932),
            .in2(N__21448),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_3_8_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_8_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_8_1  (
            .in0(_gnd_net_),
            .in1(N__20905),
            .in2(N__21544),
            .in3(N__20926),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_3_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_3_8_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_3_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_3_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20899),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49974),
            .ce(),
            .sr(N__49497));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_3_9_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_3_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJ31_LC_3_9_0  (
            .in0(_gnd_net_),
            .in1(N__20875),
            .in2(N__22013),
            .in3(N__22005),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNICOJZ0Z31 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_3_9_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_3_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI1B791_LC_3_9_1  (
            .in0(_gnd_net_),
            .in1(N__20869),
            .in2(_gnd_net_),
            .in3(N__20863),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNI1BZ0Z791 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_3_9_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_3_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNI829A1_LC_3_9_2  (
            .in0(_gnd_net_),
            .in1(N__20860),
            .in2(_gnd_net_),
            .in3(N__20842),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNI829AZ0Z1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_3_9_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_3_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CA1_LC_3_9_3  (
            .in0(_gnd_net_),
            .in1(N__21136),
            .in2(_gnd_net_),
            .in3(N__21115),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNIB8CAZ0Z1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_3_9_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_3_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFA1_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(N__21259),
            .in2(_gnd_net_),
            .in3(N__21112),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNIEEFAZ0Z1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_3_9_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_3_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAO1_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(N__21922),
            .in2(_gnd_net_),
            .in3(N__21109),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIVTAOZ0Z1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_3_9_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_3_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4TP61_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(N__21019),
            .in2(_gnd_net_),
            .in3(N__21106),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNI4TPZ0Z61 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_3_9_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_3_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI85U61_LC_3_9_7  (
            .in0(_gnd_net_),
            .in1(N__21103),
            .in2(_gnd_net_),
            .in3(N__21097),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNI85UZ0Z61 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_3_10_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_3_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICD271_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__21094),
            .in2(_gnd_net_),
            .in3(N__21088),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNICDZ0Z271 ),
            .ltout(),
            .carryin(bfn_3_10_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_3_10_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_3_10_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGL671_LC_3_10_1  (
            .in0(N__21085),
            .in1(N__21079),
            .in2(N__22015),
            .in3(N__21067),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGLZ0Z671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_10_3  (
            .in0(N__22608),
            .in1(N__22502),
            .in2(N__22579),
            .in3(N__21271),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_3_10_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_3_10_4 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNI378N_LC_3_10_4  (
            .in0(N__21064),
            .in1(N__22009),
            .in2(N__21046),
            .in3(N__21025),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_10_5 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_10_5  (
            .in0(N__22650),
            .in1(N__22524),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_3_10_6  (
            .in0(N__21840),
            .in1(N__21915),
            .in2(N__21879),
            .in3(N__21661),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_3_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_3_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_3_10_7 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNIFSVQ_LC_3_10_7  (
            .in0(N__21265),
            .in1(N__21220),
            .in2(N__22014),
            .in3(N__21205),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_0 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_3_11_0  (
            .in0(N__23165),
            .in1(N__21246),
            .in2(N__22240),
            .in3(N__22329),
            .lcout(\current_shift_inst.PI_CTRL.N_153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_11_2 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_3_11_2  (
            .in0(N__23167),
            .in1(N__22692),
            .in2(N__22230),
            .in3(N__22096),
            .lcout(\current_shift_inst.PI_CTRL.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_3_11_6  (
            .in0(N__23166),
            .in1(_gnd_net_),
            .in2(N__22231),
            .in3(N__22095),
            .lcout(\current_shift_inst.PI_CTRL.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_12_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_12_5  (
            .in0(N__21197),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21216),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_3_30_2 (
            .in0(N__21181),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_4_7_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_4_7_6 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI0UJ15_LC_4_7_6  (
            .in0(N__21600),
            .in1(N__21154),
            .in2(N__21433),
            .in3(N__21807),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_4_8_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_4_8_0 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNI4R655_LC_4_8_0  (
            .in0(N__21806),
            .in1(N__21607),
            .in2(N__21556),
            .in3(N__21423),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_4_8_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_4_8_2 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIJ3BM5_LC_4_8_2  (
            .in0(N__21802),
            .in1(N__21603),
            .in2(N__21532),
            .in3(N__21419),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_4_8_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_4_8_3 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIO2Q45_LC_4_8_3  (
            .in0(N__21604),
            .in1(N__21514),
            .in2(N__21431),
            .in3(N__21803),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_4_8_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_4_8_4 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI2KF85_LC_4_8_4  (
            .in0(N__21801),
            .in1(N__21602),
            .in2(N__21496),
            .in3(N__21418),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_4_8_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_4_8_5 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNILG775_LC_4_8_5  (
            .in0(N__21601),
            .in1(N__21478),
            .in2(N__21430),
            .in3(N__21800),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_4_8_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_4_8_6 .LUT_INIT=16'b1111010111110011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNI0J255_LC_4_8_6  (
            .in0(N__21805),
            .in1(N__21606),
            .in2(N__21463),
            .in3(N__21424),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_4_8_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_4_8_7 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNISAU45_LC_4_8_7  (
            .in0(N__21605),
            .in1(N__21439),
            .in2(N__21432),
            .in3(N__21804),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_9_0 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_4_9_0  (
            .in0(N__22189),
            .in1(N__22607),
            .in2(N__22542),
            .in3(N__22571),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_4_9_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_4_9_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIV9Q81_LC_4_9_4  (
            .in0(N__22072),
            .in1(N__22063),
            .in2(N__22036),
            .in3(N__21999),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_9_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_9_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_4_9_5  (
            .in0(N__21916),
            .in1(N__21880),
            .in2(N__21727),
            .in3(N__21844),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_9_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_9_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_4_9_6  (
            .in0(N__21691),
            .in1(N__22383),
            .in2(N__21817),
            .in3(N__21648),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_4_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_4_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_4_10_3 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_4_10_3  (
            .in0(N__22257),
            .in1(N__21761),
            .in2(N__22174),
            .in3(N__22405),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49967),
            .ce(),
            .sr(N__49506));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_4_10_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_4_10_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_4_10_5  (
            .in0(N__21723),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21686),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_4_10_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_4_10_7 .LUT_INIT=16'b1010111110101011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_4_10_7  (
            .in0(N__21655),
            .in1(N__22382),
            .in2(N__21649),
            .in3(N__21616),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_11_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(N__22777),
            .in2(_gnd_net_),
            .in3(N__22800),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_11_1  (
            .in0(N__22941),
            .in1(N__22288),
            .in2(N__21562),
            .in3(N__22918),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_4_11_2  (
            .in0(N__22300),
            .in1(N__22282),
            .in2(N__21559),
            .in3(N__22246),
            .lcout(\current_shift_inst.PI_CTRL.N_53 ),
            .ltout(\current_shift_inst.PI_CTRL.N_53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_4_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_4_11_3 .LUT_INIT=16'b0100010101000100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_4_11_3  (
            .in0(N__22725),
            .in1(N__22156),
            .in2(N__22270),
            .in3(N__22138),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_4_11_4  (
            .in0(N__23052),
            .in1(N__22447),
            .in2(N__23074),
            .in3(N__23245),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_4_11_6  (
            .in0(N__22690),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22724),
            .lcout(\current_shift_inst.PI_CTRL.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_4_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_4_11_7 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_4_11_7  (
            .in0(N__22223),
            .in1(N__23142),
            .in2(_gnd_net_),
            .in3(N__22691),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_4_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_4_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_4_13_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_4_13_2  (
            .in0(N__26207),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22207),
            .ce(),
            .sr(N__49521));
    defparam \delay_measurement_inst.start_timer_hc_LC_4_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_4_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_4_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26206),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22207),
            .ce(),
            .sr(N__49521));
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_7_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_7_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D1_LC_5_7_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH2_MAX_D1_LC_5_7_1 (
            .in0(N__22198),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49972),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_5_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_5_9_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(N__22503),
            .in2(_gnd_net_),
            .in3(N__22640),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_5_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_5_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_5_10_5 .LUT_INIT=16'b1111111101010001;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_5_10_5  (
            .in0(N__22175),
            .in1(N__22137),
            .in2(N__22118),
            .in3(N__22726),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49962),
            .ce(),
            .sr(N__49498));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_5_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_5_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_5_11_0  (
            .in0(N__23244),
            .in1(N__22306),
            .in2(N__22942),
            .in3(N__22294),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_11_1  (
            .in0(N__22276),
            .in1(N__22312),
            .in2(N__22363),
            .in3(N__22453),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_11_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_11_2  (
            .in0(N__23094),
            .in1(N__22872),
            .in2(N__22896),
            .in3(N__22746),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_5_11_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_5_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_5_11_3  (
            .in0(N__23013),
            .in1(N__23028),
            .in2(N__23221),
            .in3(N__23070),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_5_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_5_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_5_11_4  (
            .in0(N__23029),
            .in1(N__22873),
            .in2(N__22897),
            .in3(N__23014),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_5_11_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_5_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__22917),
            .in2(_gnd_net_),
            .in3(N__22470),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_11_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_5_11_7  (
            .in0(N__22471),
            .in1(N__22824),
            .in2(N__22855),
            .in3(N__23220),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_5_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_5_12_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_5_12_1  (
            .in0(N__22996),
            .in1(N__23098),
            .in2(N__22981),
            .in3(N__22750),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_5_12_2  (
            .in0(N__23194),
            .in1(N__22776),
            .in2(N__22960),
            .in3(N__22801),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_5_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_5_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_5_12_5  (
            .in0(N__22995),
            .in1(N__23053),
            .in2(N__22980),
            .in3(N__22441),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__23193),
            .in2(_gnd_net_),
            .in3(N__22959),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_5_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_5_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__22825),
            .in2(_gnd_net_),
            .in3(N__22851),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_7_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_7_6_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_7_6_7 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_7_6_7  (
            .in0(N__37664),
            .in1(N__37285),
            .in2(_gnd_net_),
            .in3(N__26689),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49970),
            .ce(),
            .sr(N__49452));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_7_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_7_8_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1HI5_22_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(N__29841),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_7_8_3  (
            .in0(N__30312),
            .in1(N__35456),
            .in2(N__33813),
            .in3(N__29714),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_7_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_7_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_7_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__25411),
            .in2(N__24577),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .clk(N__49957),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_7_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_7_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_7_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__25402),
            .in2(N__29434),
            .in3(N__22408),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(N__49957),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_7_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_7_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_7_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__29257),
            .in2(N__25423),
            .in3(N__22393),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__49957),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_7_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_7_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_7_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(N__23407),
            .in2(N__34801),
            .in3(N__22699),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__49957),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__23413),
            .in2(N__29587),
            .in3(N__22660),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__49957),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(N__23395),
            .in2(N__29641),
            .in3(N__22618),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__49957),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__23419),
            .in2(N__29347),
            .in3(N__22582),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__49957),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(N__23401),
            .in2(N__33955),
            .in3(N__22546),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__49957),
            .ce(),
            .sr(N__49474));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__25459),
            .in2(N__37114),
            .in3(N__22510),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__49951),
            .ce(),
            .sr(N__49484));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__24640),
            .in2(N__38110),
            .in3(N__22474),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__49951),
            .ce(),
            .sr(N__49484));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__24667),
            .in2(N__33871),
            .in3(N__22456),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__49951),
            .ce(),
            .sr(N__49484));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(N__24649),
            .in2(N__35284),
            .in3(N__22921),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__49951),
            .ce(),
            .sr(N__49484));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__25393),
            .in2(N__29797),
            .in3(N__22900),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__49951),
            .ce(),
            .sr(N__49484));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__24658),
            .in2(N__38179),
            .in3(N__22876),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__49951),
            .ce(),
            .sr(N__49484));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_10_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__25480),
            .in2(N__29215),
            .in3(N__22858),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__49951),
            .ce(),
            .sr(N__49484));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_10_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__29490),
            .in2(N__25518),
            .in3(N__22828),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__49951),
            .ce(),
            .sr(N__49484));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__25519),
            .in2(N__38041),
            .in3(N__22804),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__33718),
            .in2(N__25551),
            .in3(N__22780),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__25523),
            .in2(N__35130),
            .in3(N__22753),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__35655),
            .in2(N__25552),
            .in3(N__22729),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__25527),
            .in2(N__34015),
            .in3(N__23077),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__33817),
            .in2(N__25553),
            .in3(N__23056),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__25531),
            .in2(N__29857),
            .in3(N__23032),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__30003),
            .in2(N__25554),
            .in3(N__23017),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__49947),
            .ce(),
            .sr(N__49491));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__35457),
            .in2(N__25555),
            .in3(N__22999),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__49943),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__25538),
            .in2(N__30316),
            .in3(N__22984),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__49943),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__29718),
            .in2(N__25556),
            .in3(N__22963),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__49943),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__25542),
            .in2(N__34090),
            .in3(N__22945),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__49943),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__27148),
            .in2(N__25557),
            .in3(N__23224),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__49943),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__25546),
            .in2(N__27193),
            .in3(N__23197),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__49943),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(N__25384),
            .in2(N__25558),
            .in3(N__23182),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__49943),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_7_12_7  (
            .in0(N__37500),
            .in1(N__25550),
            .in2(_gnd_net_),
            .in3(N__23179),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49943),
            .ce(),
            .sr(N__49499));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30745),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_7_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_7_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24756),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_7_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_7_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25922),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30829),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27334),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_7_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_7_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24802),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_7_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_7_14_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_7_14_0  (
            .in0(N__31985),
            .in1(N__24834),
            .in2(N__27436),
            .in3(N__24813),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_7_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_7_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_7_14_1  (
            .in0(N__23890),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49931),
            .ce(N__27634),
            .sr(N__49509));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_7_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_7_14_6 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_7_14_6  (
            .in0(N__31986),
            .in1(N__26415),
            .in2(N__28000),
            .in3(N__32667),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_7_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_7_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30919),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_7_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_7_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30512),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_7_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_7_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31351),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25958),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26302),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_7_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_7_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26065),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_7_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_7_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31642),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_7_16_1  (
            .in0(N__32146),
            .in1(N__26474),
            .in2(N__32726),
            .in3(N__26438),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_7_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_7_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31048),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_16_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_16_3  (
            .in0(N__32141),
            .in1(N__31169),
            .in2(N__32725),
            .in3(N__31130),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_7_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_7_16_4 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_7_16_4  (
            .in0(N__30490),
            .in1(N__32140),
            .in2(N__32728),
            .in3(N__30513),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_7_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_7_16_5 .LUT_INIT=16'b1111010100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_7_16_5  (
            .in0(N__25826),
            .in1(N__32711),
            .in2(N__32155),
            .in3(N__25790),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_7_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_7_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27266),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_7_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_7_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_7_16_7  (
            .in0(N__32142),
            .in1(N__26376),
            .in2(N__32727),
            .in3(N__26330),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_7_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_7_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24884),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_7_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_7_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24942),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_17_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_17_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_17_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_7_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_7_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31168),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_7_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_7_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25825),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_7_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_7_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26368),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_7_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_7_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31781),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_7_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_7_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31543),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_7_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_7_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26473),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24704),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_19_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__23914),
            .in2(N__23862),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49903),
            .ce(N__27631),
            .sr(N__49528));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__23886),
            .in2(N__23835),
            .in3(N__23248),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49903),
            .ce(N__27631),
            .sr(N__49528));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__23805),
            .in2(N__23863),
            .in3(N__23275),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49903),
            .ce(N__27631),
            .sr(N__49528));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__23778),
            .in2(N__23836),
            .in3(N__23272),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49903),
            .ce(N__27631),
            .sr(N__49528));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__23751),
            .in2(N__23809),
            .in3(N__23269),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49903),
            .ce(N__27631),
            .sr(N__49528));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__24123),
            .in2(N__23782),
            .in3(N__23266),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49903),
            .ce(N__27631),
            .sr(N__49528));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__24099),
            .in2(N__23755),
            .in3(N__23263),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49903),
            .ce(N__27631),
            .sr(N__49528));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__24124),
            .in2(N__24076),
            .in3(N__23260),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49903),
            .ce(N__27631),
            .sr(N__49528));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__24042),
            .in2(N__24103),
            .in3(N__23257),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49898),
            .ce(N__27630),
            .sr(N__49533));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__24018),
            .in2(N__24075),
            .in3(N__23254),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49898),
            .ce(N__27630),
            .sr(N__49533));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(N__24043),
            .in2(N__23995),
            .in3(N__23251),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49898),
            .ce(N__27630),
            .sr(N__49533));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(N__23964),
            .in2(N__24022),
            .in3(N__23302),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49898),
            .ce(N__27630),
            .sr(N__49533));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_7_20_4  (
            .in0(_gnd_net_),
            .in1(N__23994),
            .in2(N__23940),
            .in3(N__23299),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49898),
            .ce(N__27630),
            .sr(N__49533));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__24351),
            .in2(N__23968),
            .in3(N__23296),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49898),
            .ce(N__27630),
            .sr(N__49533));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(N__24327),
            .in2(N__23941),
            .in3(N__23293),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49898),
            .ce(N__27630),
            .sr(N__49533));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(N__24352),
            .in2(N__24303),
            .in3(N__23290),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49898),
            .ce(N__27630),
            .sr(N__49533));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__24273),
            .in2(N__24331),
            .in3(N__23287),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_7_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49892),
            .ce(N__27628),
            .sr(N__49537));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__24249),
            .in2(N__24304),
            .in3(N__23284),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49892),
            .ce(N__27628),
            .sr(N__49537));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(N__24274),
            .in2(N__24226),
            .in3(N__23281),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49892),
            .ce(N__27628),
            .sr(N__49537));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_7_21_3  (
            .in0(_gnd_net_),
            .in1(N__24195),
            .in2(N__24253),
            .in3(N__23278),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49892),
            .ce(N__27628),
            .sr(N__49537));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_7_21_4  (
            .in0(_gnd_net_),
            .in1(N__24225),
            .in2(N__24171),
            .in3(N__23329),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49892),
            .ce(N__27628),
            .sr(N__49537));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(N__24144),
            .in2(N__24199),
            .in3(N__23326),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49892),
            .ce(N__27628),
            .sr(N__49537));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(N__24504),
            .in2(N__24172),
            .in3(N__23323),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49892),
            .ce(N__27628),
            .sr(N__49537));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(N__24145),
            .in2(N__24480),
            .in3(N__23320),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49892),
            .ce(N__27628),
            .sr(N__49537));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_7_22_0  (
            .in0(_gnd_net_),
            .in1(N__24450),
            .in2(N__24508),
            .in3(N__23317),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_7_22_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49885),
            .ce(N__27627),
            .sr(N__49541));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_7_22_1  (
            .in0(_gnd_net_),
            .in1(N__24426),
            .in2(N__24481),
            .in3(N__23314),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49885),
            .ce(N__27627),
            .sr(N__49541));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_7_22_2  (
            .in0(_gnd_net_),
            .in1(N__24451),
            .in2(N__24403),
            .in3(N__23311),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49885),
            .ce(N__27627),
            .sr(N__49541));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_7_22_3  (
            .in0(_gnd_net_),
            .in1(N__24379),
            .in2(N__24430),
            .in3(N__23308),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49885),
            .ce(N__27627),
            .sr(N__49541));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_7_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23305),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_5_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_5_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D1_LC_8_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D1_LC_8_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23380),
            .lcout(il_min_comp2_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49971),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_8_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_8_6_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_0_LC_8_6_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_0_LC_8_6_2  (
            .in0(N__37663),
            .in1(N__37234),
            .in2(_gnd_net_),
            .in3(N__26728),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49968),
            .ce(),
            .sr(N__49444));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI967M_13_LC_8_7_3  (
            .in0(N__38037),
            .in1(N__29204),
            .in2(N__38174),
            .in3(N__29997),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMJHC1_28_LC_8_7_4  (
            .in0(N__27147),
            .in1(N__23365),
            .in2(N__23368),
            .in3(N__34084),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_7_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI005B_30_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__25380),
            .in2(_gnd_net_),
            .in3(N__29793),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH2_MAX_D2_LC_8_8_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_8_8_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MAX_D2_LC_8_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MAX_D2_LC_8_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23359),
            .lcout(il_max_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49958),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFE9M_18_LC_8_8_1  (
            .in0(N__37488),
            .in1(N__35123),
            .in2(N__29852),
            .in3(N__35656),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_18_LC_8_8_2  (
            .in0(N__23347),
            .in1(N__23341),
            .in2(N__23335),
            .in3(N__23425),
            .lcout(\current_shift_inst.PI_CTRL.N_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_8_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_8_8_4  (
            .in0(N__37107),
            .in1(N__33936),
            .in2(N__29346),
            .in3(N__38103),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_8_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_8_8_5  (
            .in0(N__29582),
            .in1(N__34796),
            .in2(N__23332),
            .in3(N__29637),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_72_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHL6U3_29_LC_8_8_6  (
            .in0(N__33862),
            .in1(N__24607),
            .in2(N__23428),
            .in3(N__27185),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_8_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_8_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30148),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49952),
            .ce(),
            .sr(N__49467));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_8_9_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_8_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29916),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49952),
            .ce(),
            .sr(N__49467));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_8_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_8_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33231),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49952),
            .ce(),
            .sr(N__49467));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_8_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_8_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30119),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49952),
            .ce(),
            .sr(N__49467));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_8_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_8_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29886),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49952),
            .ce(),
            .sr(N__49467));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27485),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_12_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_8_12_5  (
            .in0(N__27486),
            .in1(_gnd_net_),
            .in2(N__23389),
            .in3(N__30656),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_8_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_8_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__23386),
            .in2(N__27527),
            .in3(N__27528),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_8_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_8_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__23725),
            .in2(_gnd_net_),
            .in3(N__23494),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_8_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_8_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__23491),
            .in2(_gnd_net_),
            .in3(N__23485),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_8_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_8_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__23482),
            .in2(_gnd_net_),
            .in3(N__23476),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_8_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_8_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__23473),
            .in2(_gnd_net_),
            .in3(N__23467),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_8_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_8_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__23464),
            .in2(_gnd_net_),
            .in3(N__23452),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_8_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_8_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__23449),
            .in2(_gnd_net_),
            .in3(N__23443),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_8_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_8_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__23440),
            .in2(_gnd_net_),
            .in3(N__23434),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_8_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_8_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__23686),
            .in2(_gnd_net_),
            .in3(N__23431),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_8_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_8_14_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23701),
            .in3(N__23563),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_8_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_8_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__23560),
            .in2(_gnd_net_),
            .in3(N__23554),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_8_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_8_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__23713),
            .in2(_gnd_net_),
            .in3(N__23551),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_8_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_8_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__23548),
            .in2(_gnd_net_),
            .in3(N__23542),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_8_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_8_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__23539),
            .in2(_gnd_net_),
            .in3(N__23533),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_8_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_8_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__23530),
            .in2(_gnd_net_),
            .in3(N__23524),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_8_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_8_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_8_14_7  (
            .in0(_gnd_net_),
            .in1(N__23521),
            .in2(_gnd_net_),
            .in3(N__23515),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_8_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_8_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__23512),
            .in2(_gnd_net_),
            .in3(N__23506),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_8_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_8_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__23503),
            .in2(_gnd_net_),
            .in3(N__23497),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_8_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_8_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__23641),
            .in2(_gnd_net_),
            .in3(N__23632),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_8_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_8_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__23629),
            .in2(_gnd_net_),
            .in3(N__23620),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_8_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_8_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__23617),
            .in2(_gnd_net_),
            .in3(N__23608),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_8_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_8_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__25843),
            .in2(_gnd_net_),
            .in3(N__23605),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_8_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_8_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__23602),
            .in2(_gnd_net_),
            .in3(N__23593),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_8_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_8_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__23590),
            .in2(_gnd_net_),
            .in3(N__23584),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_8_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_8_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(N__23581),
            .in2(_gnd_net_),
            .in3(N__23575),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_8_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_8_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(N__23572),
            .in2(_gnd_net_),
            .in3(N__23566),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_8_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_8_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_8_16_2  (
            .in0(_gnd_net_),
            .in1(N__23677),
            .in2(_gnd_net_),
            .in3(N__23671),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_8_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_8_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(N__23668),
            .in2(_gnd_net_),
            .in3(N__23662),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_8_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_8_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(N__23659),
            .in2(_gnd_net_),
            .in3(N__23650),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_8_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_8_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23647),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_8_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_8_16_6 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23644),
            .in3(N__32138),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_8_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_8_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_8_16_7  (
            .in0(N__30620),
            .in1(N__30749),
            .in2(_gnd_net_),
            .in3(N__30714),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_8_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_8_17_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_8_17_0  (
            .in0(N__30619),
            .in1(N__25995),
            .in2(_gnd_net_),
            .in3(N__25952),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_8_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_8_17_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_8_17_1  (
            .in0(N__27335),
            .in1(N__30616),
            .in2(_gnd_net_),
            .in3(N__27303),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_8_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_8_17_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_8_17_2  (
            .in0(N__32108),
            .in1(N__27267),
            .in2(_gnd_net_),
            .in3(N__27225),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_17_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_8_17_3  (
            .in0(N__25871),
            .in1(N__30618),
            .in2(_gnd_net_),
            .in3(N__25915),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_8_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_8_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_8_17_4  (
            .in0(N__30615),
            .in1(N__30830),
            .in2(_gnd_net_),
            .in3(N__30798),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_8_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_8_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_8_17_5  (
            .in0(N__30622),
            .in1(N__31406),
            .in2(_gnd_net_),
            .in3(N__31449),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_8_17_6  (
            .in0(N__30617),
            .in1(N__24711),
            .in2(_gnd_net_),
            .in3(N__24687),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_8_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_8_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_8_17_7  (
            .in0(N__30621),
            .in1(N__24752),
            .in2(_gnd_net_),
            .in3(N__24787),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_8_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_8_18_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_8_18_0  (
            .in0(N__30923),
            .in1(N__30643),
            .in2(_gnd_net_),
            .in3(N__30888),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_8_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_8_18_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_8_18_1  (
            .in0(N__30645),
            .in1(N__31059),
            .in2(_gnd_net_),
            .in3(N__31088),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_8_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_8_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30981),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_8_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_8_18_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_8_18_3  (
            .in0(N__30647),
            .in1(_gnd_net_),
            .in2(N__31788),
            .in3(N__31829),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_8_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_8_18_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_8_18_4  (
            .in0(N__26066),
            .in1(N__30646),
            .in2(_gnd_net_),
            .in3(N__26028),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_8_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_8_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_8_18_5  (
            .in0(N__30648),
            .in1(N__31228),
            .in2(_gnd_net_),
            .in3(N__31266),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_8_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_8_18_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_8_18_6  (
            .in0(N__27558),
            .in1(N__30642),
            .in2(_gnd_net_),
            .in3(N__27599),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_8_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_8_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_8_18_7  (
            .in0(N__30644),
            .in1(N__26303),
            .in2(_gnd_net_),
            .in3(N__26258),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_8_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_8_19_0 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_8_19_0  (
            .in0(N__31653),
            .in1(N__31595),
            .in2(_gnd_net_),
            .in3(N__30655),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_8_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_8_19_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__27557),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_8_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_8_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26112),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_8_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_8_19_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_8_19_3  (
            .in0(N__30654),
            .in1(N__31544),
            .in2(_gnd_net_),
            .in3(N__31512),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_8_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_8_19_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_8_19_4  (
            .in0(N__32156),
            .in1(N__26369),
            .in2(_gnd_net_),
            .in3(N__26337),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_8_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_8_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31396),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_8_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_8_19_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_8_19_6  (
            .in0(N__32158),
            .in1(_gnd_net_),
            .in2(N__26481),
            .in3(N__26442),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_8_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_8_19_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_8_19_7  (
            .in0(N__25827),
            .in1(N__32157),
            .in2(_gnd_net_),
            .in3(N__25794),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23913),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49893),
            .ce(N__27629),
            .sr(N__49529));
    defparam \current_shift_inst.timer_s1.counter_0_LC_8_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_8_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_8_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_8_21_0  (
            .in0(N__25325),
            .in1(N__23912),
            .in2(_gnd_net_),
            .in3(N__23893),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__49886),
            .ce(N__33358),
            .sr(N__49534));
    defparam \current_shift_inst.timer_s1.counter_1_LC_8_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_8_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_8_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_8_21_1  (
            .in0(N__25342),
            .in1(N__23885),
            .in2(_gnd_net_),
            .in3(N__23866),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__49886),
            .ce(N__33358),
            .sr(N__49534));
    defparam \current_shift_inst.timer_s1.counter_2_LC_8_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_8_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_8_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_8_21_2  (
            .in0(N__25326),
            .in1(N__23855),
            .in2(_gnd_net_),
            .in3(N__23839),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__49886),
            .ce(N__33358),
            .sr(N__49534));
    defparam \current_shift_inst.timer_s1.counter_3_LC_8_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_8_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_8_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_8_21_3  (
            .in0(N__25343),
            .in1(N__23828),
            .in2(_gnd_net_),
            .in3(N__23812),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__49886),
            .ce(N__33358),
            .sr(N__49534));
    defparam \current_shift_inst.timer_s1.counter_4_LC_8_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_8_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_8_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_8_21_4  (
            .in0(N__25327),
            .in1(N__23804),
            .in2(_gnd_net_),
            .in3(N__23785),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__49886),
            .ce(N__33358),
            .sr(N__49534));
    defparam \current_shift_inst.timer_s1.counter_5_LC_8_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_8_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_8_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_8_21_5  (
            .in0(N__25344),
            .in1(N__23777),
            .in2(_gnd_net_),
            .in3(N__23758),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__49886),
            .ce(N__33358),
            .sr(N__49534));
    defparam \current_shift_inst.timer_s1.counter_6_LC_8_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_8_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_8_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_8_21_6  (
            .in0(N__25328),
            .in1(N__23744),
            .in2(_gnd_net_),
            .in3(N__23728),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__49886),
            .ce(N__33358),
            .sr(N__49534));
    defparam \current_shift_inst.timer_s1.counter_7_LC_8_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_8_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_8_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_8_21_7  (
            .in0(N__25345),
            .in1(N__24122),
            .in2(_gnd_net_),
            .in3(N__24106),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__49886),
            .ce(N__33358),
            .sr(N__49534));
    defparam \current_shift_inst.timer_s1.counter_8_LC_8_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_8_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_8_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_8_22_0  (
            .in0(N__25324),
            .in1(N__24098),
            .in2(_gnd_net_),
            .in3(N__24079),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__49879),
            .ce(N__33356),
            .sr(N__49538));
    defparam \current_shift_inst.timer_s1.counter_9_LC_8_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_8_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_8_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_8_22_1  (
            .in0(N__25332),
            .in1(N__24065),
            .in2(_gnd_net_),
            .in3(N__24046),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__49879),
            .ce(N__33356),
            .sr(N__49538));
    defparam \current_shift_inst.timer_s1.counter_10_LC_8_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_8_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_8_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_8_22_2  (
            .in0(N__25321),
            .in1(N__24041),
            .in2(_gnd_net_),
            .in3(N__24025),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__49879),
            .ce(N__33356),
            .sr(N__49538));
    defparam \current_shift_inst.timer_s1.counter_11_LC_8_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_8_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_8_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_8_22_3  (
            .in0(N__25329),
            .in1(N__24017),
            .in2(_gnd_net_),
            .in3(N__23998),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__49879),
            .ce(N__33356),
            .sr(N__49538));
    defparam \current_shift_inst.timer_s1.counter_12_LC_8_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_8_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_8_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_8_22_4  (
            .in0(N__25322),
            .in1(N__23990),
            .in2(_gnd_net_),
            .in3(N__23971),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__49879),
            .ce(N__33356),
            .sr(N__49538));
    defparam \current_shift_inst.timer_s1.counter_13_LC_8_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_8_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_8_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_8_22_5  (
            .in0(N__25330),
            .in1(N__23963),
            .in2(_gnd_net_),
            .in3(N__23944),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__49879),
            .ce(N__33356),
            .sr(N__49538));
    defparam \current_shift_inst.timer_s1.counter_14_LC_8_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_8_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_8_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_8_22_6  (
            .in0(N__25323),
            .in1(N__23933),
            .in2(_gnd_net_),
            .in3(N__23917),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__49879),
            .ce(N__33356),
            .sr(N__49538));
    defparam \current_shift_inst.timer_s1.counter_15_LC_8_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_8_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_8_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_8_22_7  (
            .in0(N__25331),
            .in1(N__24350),
            .in2(_gnd_net_),
            .in3(N__24334),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__49879),
            .ce(N__33356),
            .sr(N__49538));
    defparam \current_shift_inst.timer_s1.counter_16_LC_8_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_8_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_8_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_8_23_0  (
            .in0(N__25311),
            .in1(N__24326),
            .in2(_gnd_net_),
            .in3(N__24307),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_23_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__49871),
            .ce(N__33357),
            .sr(N__49542));
    defparam \current_shift_inst.timer_s1.counter_17_LC_8_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_8_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_8_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_8_23_1  (
            .in0(N__25315),
            .in1(N__24296),
            .in2(_gnd_net_),
            .in3(N__24277),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__49871),
            .ce(N__33357),
            .sr(N__49542));
    defparam \current_shift_inst.timer_s1.counter_18_LC_8_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_8_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_8_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_8_23_2  (
            .in0(N__25312),
            .in1(N__24272),
            .in2(_gnd_net_),
            .in3(N__24256),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__49871),
            .ce(N__33357),
            .sr(N__49542));
    defparam \current_shift_inst.timer_s1.counter_19_LC_8_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_8_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_8_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_8_23_3  (
            .in0(N__25316),
            .in1(N__24248),
            .in2(_gnd_net_),
            .in3(N__24229),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__49871),
            .ce(N__33357),
            .sr(N__49542));
    defparam \current_shift_inst.timer_s1.counter_20_LC_8_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_8_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_8_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_8_23_4  (
            .in0(N__25313),
            .in1(N__24221),
            .in2(_gnd_net_),
            .in3(N__24202),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__49871),
            .ce(N__33357),
            .sr(N__49542));
    defparam \current_shift_inst.timer_s1.counter_21_LC_8_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_8_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_8_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_8_23_5  (
            .in0(N__25317),
            .in1(N__24194),
            .in2(_gnd_net_),
            .in3(N__24175),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__49871),
            .ce(N__33357),
            .sr(N__49542));
    defparam \current_shift_inst.timer_s1.counter_22_LC_8_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_8_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_8_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_8_23_6  (
            .in0(N__25314),
            .in1(N__24164),
            .in2(_gnd_net_),
            .in3(N__24148),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__49871),
            .ce(N__33357),
            .sr(N__49542));
    defparam \current_shift_inst.timer_s1.counter_23_LC_8_23_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_8_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_8_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_8_23_7  (
            .in0(N__25318),
            .in1(N__24143),
            .in2(_gnd_net_),
            .in3(N__24127),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__49871),
            .ce(N__33357),
            .sr(N__49542));
    defparam \current_shift_inst.timer_s1.counter_24_LC_8_24_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_8_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_8_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_8_24_0  (
            .in0(N__25307),
            .in1(N__24503),
            .in2(_gnd_net_),
            .in3(N__24484),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_24_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__49867),
            .ce(N__33341),
            .sr(N__49543));
    defparam \current_shift_inst.timer_s1.counter_25_LC_8_24_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_8_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_8_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_8_24_1  (
            .in0(N__25319),
            .in1(N__24473),
            .in2(_gnd_net_),
            .in3(N__24454),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__49867),
            .ce(N__33341),
            .sr(N__49543));
    defparam \current_shift_inst.timer_s1.counter_26_LC_8_24_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_8_24_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_8_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_8_24_2  (
            .in0(N__25308),
            .in1(N__24449),
            .in2(_gnd_net_),
            .in3(N__24433),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__49867),
            .ce(N__33341),
            .sr(N__49543));
    defparam \current_shift_inst.timer_s1.counter_27_LC_8_24_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_8_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_8_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_8_24_3  (
            .in0(N__25320),
            .in1(N__24425),
            .in2(_gnd_net_),
            .in3(N__24406),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__49867),
            .ce(N__33341),
            .sr(N__49543));
    defparam \current_shift_inst.timer_s1.counter_28_LC_8_24_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_8_24_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_8_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_8_24_4  (
            .in0(N__25309),
            .in1(N__24399),
            .in2(_gnd_net_),
            .in3(N__24385),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__49867),
            .ce(N__33341),
            .sr(N__49543));
    defparam \current_shift_inst.timer_s1.counter_29_LC_8_24_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_8_24_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_8_24_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_8_24_5  (
            .in0(N__24375),
            .in1(N__25310),
            .in2(_gnd_net_),
            .in3(N__24382),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49867),
            .ce(N__33341),
            .sr(N__49543));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_5_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJF8D_6_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29338),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_5_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_5_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_9_5_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_9_5_4 (
            .in0(N__24361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49969),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_9_5_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_9_5_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAVO71_0_LC_9_5_5  (
            .in0(N__29262),
            .in1(N__29416),
            .in2(_gnd_net_),
            .in3(N__24570),
            .lcout(\current_shift_inst.PI_CTRL.un1_enablelt3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_9_5_6.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_9_5_6.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_9_5_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_9_5_6 (
            .in0(N__24589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49969),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_9_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_9_6_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIC35V7_13_LC_9_6_0  (
            .in0(N__24553),
            .in1(N__24613),
            .in2(N__24520),
            .in3(N__24541),
            .lcout(\current_shift_inst.PI_CTRL.N_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_6_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID98D_0_LC_9_6_2  (
            .in0(N__24569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_9_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_9_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI967M_0_13_LC_9_6_3  (
            .in0(N__38036),
            .in1(N__29203),
            .in2(N__38178),
            .in3(N__29998),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_9_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_9_6_5 .LUT_INIT=16'b1111010011110101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFCK44_3_LC_9_6_5  (
            .in0(N__29566),
            .in1(N__24547),
            .in2(N__24532),
            .in3(N__34797),
            .lcout(\current_shift_inst.PI_CTRL.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_6_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6VGQ_5_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__33950),
            .in2(_gnd_net_),
            .in3(N__29633),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_6_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JA22_6_LC_9_6_7  (
            .in0(N__38095),
            .in1(N__37100),
            .in2(N__24535),
            .in3(N__29328),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_9_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_9_7_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI654B_29_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__27175),
            .in2(_gnd_net_),
            .in3(N__33863),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_9_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_9_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID8UD2_11_LC_9_7_1  (
            .in0(N__24601),
            .in1(N__24619),
            .in2(N__24523),
            .in3(N__24595),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0FH5_12_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29784),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_9_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_9_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHF8M_18_LC_9_7_6  (
            .in0(N__35446),
            .in1(N__35634),
            .in2(N__29842),
            .in3(N__35104),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_9_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_9_7_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI78BM_30_LC_9_7_7  (
            .in0(N__34085),
            .in1(N__29785),
            .in2(N__25379),
            .in3(N__37444),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_9_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_9_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_11_LC_9_8_0  (
            .in0(N__33703),
            .in1(N__35265),
            .in2(N__29482),
            .in3(N__34006),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_9_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_9_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGGAM_28_LC_9_8_2  (
            .in0(N__27133),
            .in1(N__30304),
            .in2(N__33812),
            .in3(N__29703),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6MI5_27_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34060),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI637M_0_11_LC_9_8_4  (
            .in0(N__33702),
            .in1(N__35266),
            .in2(N__29483),
            .in3(N__34007),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI6LH5_18_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35103),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_9_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_9_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0HJ5_30_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25375),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_9_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_9_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIKG8D_7_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33949),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_9_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_9_9_6 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_9_9_6  (
            .in0(N__37439),
            .in1(N__37283),
            .in2(N__37665),
            .in3(N__27046),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49948),
            .ce(),
            .sr(N__49461));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_9_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_9_9_7 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_9_9_7  (
            .in0(N__37282),
            .in1(N__37440),
            .in2(N__27034),
            .in3(N__37602),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49948),
            .ce(),
            .sr(N__49461));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_9_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_9_10_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__30058),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49944),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_9_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_9_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33753),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49944),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_9_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_9_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30034),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49944),
            .ce(),
            .sr(N__49468));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_9_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_9_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35018),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49944),
            .ce(),
            .sr(N__49468));
    defparam SB_DFF_inst_PH2_MIN_D2_LC_9_12_4.C_ON=1'b0;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_9_12_4.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH2_MIN_D2_LC_9_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH2_MIN_D2_LC_9_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24631),
            .lcout(il_min_comp2_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49932),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32853),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_9_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_9_13_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_9_13_0  (
            .in0(N__32642),
            .in1(N__32090),
            .in2(N__24724),
            .in3(N__24683),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_9_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_9_13_1 .LUT_INIT=16'b1100010111000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_9_13_1  (
            .in0(N__24763),
            .in1(N__24782),
            .in2(N__32139),
            .in3(N__32645),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_9_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_9_13_2 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_9_13_2  (
            .in0(N__32644),
            .in1(N__32092),
            .in2(N__24786),
            .in3(N__24762),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_9_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_9_13_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_9_13_3  (
            .in0(N__32088),
            .in1(N__32640),
            .in2(N__27352),
            .in3(N__27299),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_9_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_9_13_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_9_13_4  (
            .in0(N__32641),
            .in1(N__32089),
            .in2(N__30765),
            .in3(N__30713),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_13_5 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_9_13_5  (
            .in0(N__32086),
            .in1(N__27432),
            .in2(N__24838),
            .in3(N__24817),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_9_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_9_13_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_9_13_6  (
            .in0(N__32639),
            .in1(N__32087),
            .in2(N__30850),
            .in3(N__30791),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_9_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_9_13_7 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_9_13_7  (
            .in0(N__32091),
            .in1(N__24723),
            .in2(N__24688),
            .in3(N__32643),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_9_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_9_14_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_9_14_0  (
            .in0(N__32717),
            .in1(N__31990),
            .in2(N__30535),
            .in3(N__30485),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_9_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_9_14_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_9_14_1  (
            .in0(N__31992),
            .in1(N__32719),
            .in2(N__30939),
            .in3(N__30884),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_14_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_9_14_2  (
            .in0(N__30657),
            .in1(N__24833),
            .in2(_gnd_net_),
            .in3(N__24812),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_9_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_9_14_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_9_14_3  (
            .in0(N__31987),
            .in1(N__32721),
            .in2(N__25879),
            .in3(N__25923),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_9_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_9_14_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_9_14_4  (
            .in0(N__32720),
            .in1(N__31993),
            .in2(N__31369),
            .in3(N__31301),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_9_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_9_14_5 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_9_14_5  (
            .in0(N__31988),
            .in1(N__30963),
            .in2(N__31014),
            .in3(N__32722),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_9_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_9_14_6 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_9_14_6  (
            .in0(N__32716),
            .in1(N__31442),
            .in2(N__31423),
            .in3(N__31989),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_9_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_9_14_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_9_14_7  (
            .in0(N__31991),
            .in1(N__32718),
            .in2(N__26137),
            .in3(N__26094),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_9_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_9_15_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_9_15_0  (
            .in0(N__32114),
            .in1(N__32637),
            .in2(N__25971),
            .in3(N__25994),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_15_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_9_15_1  (
            .in0(N__26133),
            .in1(N__30624),
            .in2(_gnd_net_),
            .in3(N__26093),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_9_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_9_15_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_9_15_2  (
            .in0(N__32117),
            .in1(N__32634),
            .in2(N__31243),
            .in3(N__31262),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_9_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_9_15_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_9_15_3  (
            .in0(N__32635),
            .in1(N__32118),
            .in2(N__31564),
            .in3(N__31508),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_9_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_9_15_4 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_9_15_4  (
            .in0(N__32119),
            .in1(N__31652),
            .in2(N__31612),
            .in3(N__32636),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_9_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_9_15_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_9_15_5  (
            .in0(N__32638),
            .in1(N__32115),
            .in2(N__26077),
            .in3(N__26021),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_15_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_9_15_6  (
            .in0(N__30623),
            .in1(N__31001),
            .in2(_gnd_net_),
            .in3(N__30962),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_9_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_9_15_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_9_15_7  (
            .in0(N__32633),
            .in1(N__32116),
            .in2(N__24904),
            .in3(N__24858),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_16_0 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_9_16_0  (
            .in0(N__32122),
            .in1(N__24954),
            .in2(N__24925),
            .in3(N__32673),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_9_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_9_16_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_9_16_1  (
            .in0(N__24955),
            .in1(N__24921),
            .in2(N__32715),
            .in3(N__32123),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_9_16_2  (
            .in0(N__32120),
            .in1(N__24953),
            .in2(_gnd_net_),
            .in3(N__24915),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_9_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_9_16_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_9_16_3  (
            .in0(N__32672),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32124),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_16_4 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_9_16_4  (
            .in0(N__32121),
            .in1(N__32677),
            .in2(N__24859),
            .in3(N__24900),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_16_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_9_16_6  (
            .in0(N__30630),
            .in1(N__24899),
            .in2(_gnd_net_),
            .in3(N__24854),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_9_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_9_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_9_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27666),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49909),
            .ce(N__27633),
            .sr(N__49510));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_9_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__27995),
            .in2(N__26541),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_9_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(N__28070),
            .in2(N__25012),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_9_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(N__25000),
            .in2(N__28164),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_9_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(N__28074),
            .in2(N__24994),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_9_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_9_17_4  (
            .in0(_gnd_net_),
            .in1(N__24985),
            .in2(N__28165),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_9_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(N__28078),
            .in2(N__24979),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_9_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(N__24970),
            .in2(N__28166),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_9_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(N__28082),
            .in2(N__24964),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_9_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__28179),
            .in2(N__25066),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_9_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__25057),
            .in2(N__28269),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_9_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__28167),
            .in2(N__25048),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_9_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__30463),
            .in2(N__28266),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_9_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__28171),
            .in2(N__25036),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_9_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__25024),
            .in2(N__28267),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_9_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__28175),
            .in2(N__26389),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_9_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__25018),
            .in2(N__28268),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_9_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__28183),
            .in2(N__25120),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_9_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__25111),
            .in2(N__28270),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_9_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__28187),
            .in2(N__25105),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_9_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__25096),
            .in2(N__28271),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_9_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__28191),
            .in2(N__26398),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_9_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__25090),
            .in2(N__28272),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_9_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__28195),
            .in2(N__25081),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_9_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__25072),
            .in2(N__28273),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_9_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__28199),
            .in2(N__25204),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_9_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__25195),
            .in2(N__28274),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_9_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__28203),
            .in2(N__25189),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_9_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__25180),
            .in2(N__28275),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_9_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__28207),
            .in2(N__25171),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_9_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__25156),
            .in2(N__28276),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_9_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__28211),
            .in2(N__25150),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__32147),
            .in2(_gnd_net_),
            .in3(N__25135),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S1_LC_9_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41261),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49880),
            .ce(),
            .sr(N__49530));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34879),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_9_28_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_9_28_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_9_28_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_9_28_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35884),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49851),
            .ce(),
            .sr(N__49544));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_4_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_4_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_10_4_1 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_10_4_1  (
            .in0(N__37673),
            .in1(N__37307),
            .in2(_gnd_net_),
            .in3(N__26707),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49963),
            .ce(),
            .sr(N__49414));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_5_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_5_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_10_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25210),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49959),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEA8D_1_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29420),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_10_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_10_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2HH5_14_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29193),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_10_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_10_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3IH5_15_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29481),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIFB8D_2_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29261),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHD8D_4_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29559),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_10_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_10_7_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_10_7_2 .LUT_INIT=16'b0000110011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_10_7_2  (
            .in0(N__37230),
            .in1(N__37456),
            .in2(N__37706),
            .in3(N__26647),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49949),
            .ce(),
            .sr(N__49430));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_10_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_10_7_3 .LUT_INIT=16'b0000111110101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_10_7_3  (
            .in0(N__37453),
            .in1(N__37231),
            .in2(N__26743),
            .in3(N__37686),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49949),
            .ce(),
            .sr(N__49430));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_7_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_7_5 .LUT_INIT=16'b0000111110101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_10_7_5  (
            .in0(N__37454),
            .in1(N__37232),
            .in2(N__26926),
            .in3(N__37687),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49949),
            .ce(),
            .sr(N__49430));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_10_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_10_7_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_10_7_7 .LUT_INIT=16'b0000111110101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_10_7_7  (
            .in0(N__37455),
            .in1(N__37233),
            .in2(N__26857),
            .in3(N__37688),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49949),
            .ce(),
            .sr(N__49430));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_8_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_8_0 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_10_8_0  (
            .in0(N__37269),
            .in1(N__37452),
            .in2(N__26947),
            .in3(N__37629),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(),
            .sr(N__49437));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_10_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_10_8_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_10_8_1 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_10_8_1  (
            .in0(N__37447),
            .in1(N__37272),
            .in2(N__37671),
            .in3(N__26980),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(),
            .sr(N__49437));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_10_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_10_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_10_8_2 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_10_8_2  (
            .in0(N__37267),
            .in1(N__37450),
            .in2(N__26869),
            .in3(N__37628),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(),
            .sr(N__49437));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_10_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_10_8_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_10_8_3 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_10_8_3  (
            .in0(N__37445),
            .in1(N__37270),
            .in2(N__37669),
            .in3(N__26761),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(),
            .sr(N__49437));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_10_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_10_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_10_8_4 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_10_8_4  (
            .in0(N__37266),
            .in1(N__37449),
            .in2(N__26905),
            .in3(N__37627),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(),
            .sr(N__49437));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_10_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_10_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_10_8_5 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_10_8_5  (
            .in0(N__37448),
            .in1(N__37273),
            .in2(N__37672),
            .in3(N__26971),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(),
            .sr(N__49437));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_10_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_10_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_10_8_6 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_10_8_6  (
            .in0(N__37268),
            .in1(N__37451),
            .in2(N__26827),
            .in3(N__37630),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(),
            .sr(N__49437));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_10_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_10_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_10_8_7 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_10_8_7  (
            .in0(N__37446),
            .in1(N__37271),
            .in2(N__37670),
            .in3(N__26890),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49945),
            .ce(),
            .sr(N__49437));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_10_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_10_9_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_10_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33258),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49448));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_10_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_10_9_3 .LUT_INIT=16'b0101111101010100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_10_9_3  (
            .in0(N__26989),
            .in1(N__37308),
            .in2(N__37708),
            .in3(N__37442),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49448));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_10_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_10_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_10_9_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_10_9_4  (
            .in0(N__33312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49448));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_9_5 .LUT_INIT=16'b0100010001010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_10_9_5  (
            .in0(N__26806),
            .in1(N__37693),
            .in2(N__37325),
            .in3(N__37443),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49448));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_10_9_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_10_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_10_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33288),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49448));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_10_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_10_9_7 .LUT_INIT=16'b0111011101010100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_10_9_7  (
            .in0(N__27016),
            .in1(N__37692),
            .in2(N__37324),
            .in3(N__37441),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49937),
            .ce(),
            .sr(N__49448));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_10_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_10_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_10_10_1  (
            .in0(N__35183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49933),
            .ce(),
            .sr(N__49456));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_10_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_10_10_3 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_10_10_3  (
            .in0(N__37315),
            .in1(N__37438),
            .in2(N__27202),
            .in3(N__37682),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49933),
            .ce(),
            .sr(N__49456));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_10_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_10_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37932),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49933),
            .ce(),
            .sr(N__49456));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_10_10_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_10_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_10_10_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__30090),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49933),
            .ce(),
            .sr(N__49456));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_10_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_10_12_4 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_10_12_4  (
            .in0(N__28998),
            .in1(N__35366),
            .in2(_gnd_net_),
            .in3(N__29059),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49919),
            .ce(),
            .sr(N__49469));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_10_12_6 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_10_12_6  (
            .in0(N__32881),
            .in1(N__26223),
            .in2(_gnd_net_),
            .in3(N__26185),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49919),
            .ce(),
            .sr(N__49469));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_10_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_10_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__27925),
            .in2(N__27942),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_10_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_10_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__27422),
            .in2(N__25447),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_10_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_10_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__32598),
            .in2(N__27541),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_10_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_10_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__25438),
            .in2(N__32669),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_10_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_10_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__32602),
            .in2(N__25432),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_10_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_10_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__25624),
            .in2(N__32670),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_10_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_10_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__32606),
            .in2(N__25618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_10_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_10_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__25609),
            .in2(N__32671),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_10_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_10_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__32330),
            .in2(N__25603),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_10_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_10_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__25594),
            .in2(N__32525),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_10_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_10_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__32334),
            .in2(N__25588),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_10_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_10_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__25579),
            .in2(N__32526),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_10_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_10_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__32338),
            .in2(N__25573),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_10_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_10_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__25564),
            .in2(N__32527),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_10_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_10_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__32342),
            .in2(N__25660),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_10_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_10_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__25651),
            .in2(N__32528),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_10_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_10_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__32362),
            .in2(N__26236),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_10_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_10_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__31024),
            .in2(N__32533),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_10_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_10_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__32366),
            .in2(N__25645),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_10_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_10_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__30859),
            .in2(N__32534),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_10_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_10_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__32370),
            .in2(N__31111),
            .in3(N__25636),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_10_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_10_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__25633),
            .in2(N__32535),
            .in3(N__25627),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_10_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_10_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__32374),
            .in2(N__25771),
            .in3(N__25759),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_10_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_10_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__25756),
            .in2(N__32536),
            .in3(N__25750),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_10_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_10_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__32431),
            .in2(N__25747),
            .in3(N__25738),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_10_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_10_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__25735),
            .in2(N__32585),
            .in3(N__25726),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_10_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_10_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__32435),
            .in2(N__25723),
            .in3(N__25711),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_10_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_10_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__27214),
            .in2(N__32586),
            .in3(N__25708),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_10_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_10_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__32439),
            .in2(N__25705),
            .in3(N__25693),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_10_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_10_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__25690),
            .in2(N__32587),
            .in3(N__25681),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_10_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_10_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__32443),
            .in2(N__25678),
            .in3(N__25663),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_10_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_10_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_10_16_7  (
            .in0(N__32444),
            .in1(N__32128),
            .in2(_gnd_net_),
            .in3(N__26140),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_10_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_10_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_10_17_0  (
            .in0(N__32015),
            .in1(N__26132),
            .in2(N__32653),
            .in3(N__26101),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_10_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_10_17_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_10_17_1  (
            .in0(N__31063),
            .in1(N__32018),
            .in2(N__31099),
            .in3(N__32571),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_10_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_10_17_3 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_10_17_3  (
            .in0(N__26310),
            .in1(N__32017),
            .in2(N__26272),
            .in3(N__32570),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_10_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_10_17_4 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_10_17_4  (
            .in0(N__32572),
            .in1(N__26076),
            .in2(N__32107),
            .in3(N__26032),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_17_5 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_10_17_5  (
            .in0(N__25999),
            .in1(N__32569),
            .in2(N__25975),
            .in3(N__32016),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_10_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_10_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_10_17_6  (
            .in0(N__32014),
            .in1(N__25924),
            .in2(N__32654),
            .in3(N__25875),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31232),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_18_0  (
            .in0(N__25831),
            .in1(N__32111),
            .in2(N__32724),
            .in3(N__25798),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_18_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_10_18_2  (
            .in0(N__32693),
            .in1(N__32112),
            .in2(N__26488),
            .in3(N__26446),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_10_18_3  (
            .in0(N__32113),
            .in1(N__32701),
            .in2(N__27996),
            .in3(N__26419),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_18_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_10_18_4  (
            .in0(N__31182),
            .in1(N__30653),
            .in2(_gnd_net_),
            .in3(N__31137),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_18_5  (
            .in0(N__30652),
            .in1(N__31352),
            .in2(_gnd_net_),
            .in3(N__31311),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_6  (
            .in0(N__26377),
            .in1(N__32110),
            .in2(N__32723),
            .in3(N__26341),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_10_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_10_18_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_10_18_7  (
            .in0(N__32109),
            .in1(N__32700),
            .in2(N__26314),
            .in3(N__26265),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_19_0 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_19_0  (
            .in0(N__32892),
            .in1(N__26224),
            .in2(_gnd_net_),
            .in3(N__26181),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_398_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_10_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_10_19_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__36228),
            .in2(_gnd_net_),
            .in3(N__36181),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_10_20_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_10_20_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__32891),
            .in2(_gnd_net_),
            .in3(N__26180),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_397_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_10_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_10_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_10_20_6  (
            .in0(N__26542),
            .in1(N__28212),
            .in2(_gnd_net_),
            .in3(N__26512),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27659),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49868),
            .ce(N__27626),
            .sr(N__49524));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__28927),
            .in2(N__28720),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_10_22_1  (
            .in0(N__43124),
            .in1(N__27891),
            .in2(_gnd_net_),
            .in3(N__26506),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49526));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_22_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_10_22_2  (
            .in0(N__43121),
            .in1(N__28578),
            .in2(N__28744),
            .in3(N__26503),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49526));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_10_22_3  (
            .in0(N__43125),
            .in1(N__28554),
            .in2(_gnd_net_),
            .in3(N__26500),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49526));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_10_22_4  (
            .in0(N__43122),
            .in1(N__28533),
            .in2(_gnd_net_),
            .in3(N__26497),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49526));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_10_22_5  (
            .in0(N__43126),
            .in1(N__28506),
            .in2(_gnd_net_),
            .in3(N__26494),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49526));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_10_22_6  (
            .in0(N__43123),
            .in1(N__28482),
            .in2(_gnd_net_),
            .in3(N__26491),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49526));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_22_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_10_22_7  (
            .in0(N__43127),
            .in1(N__28461),
            .in2(_gnd_net_),
            .in3(N__26569),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49863),
            .ce(),
            .sr(N__49526));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_23_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_10_23_0  (
            .in0(N__43096),
            .in1(N__28434),
            .in2(_gnd_net_),
            .in3(N__26566),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49858),
            .ce(),
            .sr(N__49531));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_10_23_1  (
            .in0(N__43089),
            .in1(N__28410),
            .in2(_gnd_net_),
            .in3(N__26563),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49858),
            .ce(),
            .sr(N__49531));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_23_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_23_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_10_23_2  (
            .in0(N__43093),
            .in1(N__28695),
            .in2(_gnd_net_),
            .in3(N__26560),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49858),
            .ce(),
            .sr(N__49531));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_23_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_10_23_3  (
            .in0(N__43090),
            .in1(N__28671),
            .in2(_gnd_net_),
            .in3(N__26557),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49858),
            .ce(),
            .sr(N__49531));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_23_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_23_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_10_23_4  (
            .in0(N__43094),
            .in1(N__28647),
            .in2(_gnd_net_),
            .in3(N__26554),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49858),
            .ce(),
            .sr(N__49531));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_10_23_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_10_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_10_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_10_23_5  (
            .in0(N__43091),
            .in1(N__28623),
            .in2(_gnd_net_),
            .in3(N__26551),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49858),
            .ce(),
            .sr(N__49531));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_23_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_10_23_6  (
            .in0(N__43095),
            .in1(N__28599),
            .in2(_gnd_net_),
            .in3(N__26548),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49858),
            .ce(),
            .sr(N__49531));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_23_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_10_23_7  (
            .in0(N__43092),
            .in1(N__42708),
            .in2(_gnd_net_),
            .in3(N__26545),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49858),
            .ce(),
            .sr(N__49531));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_24_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_24_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_10_24_0  (
            .in0(N__43139),
            .in1(N__42675),
            .in2(_gnd_net_),
            .in3(N__26596),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49535));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_24_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_24_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_10_24_1  (
            .in0(N__43132),
            .in1(N__42842),
            .in2(_gnd_net_),
            .in3(N__26593),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49535));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_24_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_24_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_10_24_2  (
            .in0(N__43140),
            .in1(N__42870),
            .in2(_gnd_net_),
            .in3(N__26590),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49535));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_10_24_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_10_24_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_10_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_10_24_3  (
            .in0(N__43133),
            .in1(N__28870),
            .in2(_gnd_net_),
            .in3(N__26587),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49535));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_10_24_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_10_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_10_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_10_24_4  (
            .in0(N__43141),
            .in1(N__28882),
            .in2(_gnd_net_),
            .in3(N__26584),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49535));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_10_24_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_10_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_10_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_10_24_5  (
            .in0(N__43134),
            .in1(N__28837),
            .in2(_gnd_net_),
            .in3(N__26581),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49535));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_10_24_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_10_24_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_10_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_10_24_6  (
            .in0(N__43142),
            .in1(N__28849),
            .in2(_gnd_net_),
            .in3(N__26578),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49535));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_10_24_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_10_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_10_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_10_24_7  (
            .in0(N__43135),
            .in1(N__28804),
            .in2(_gnd_net_),
            .in3(N__26575),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49855),
            .ce(),
            .sr(N__49535));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_10_25_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_10_25_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_10_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_10_25_0  (
            .in0(N__43128),
            .in1(N__28816),
            .in2(_gnd_net_),
            .in3(N__26572),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_10_25_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49852),
            .ce(),
            .sr(N__49539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_10_25_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_10_25_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_10_25_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_10_25_1  (
            .in0(N__43136),
            .in1(N__28771),
            .in2(_gnd_net_),
            .in3(N__26614),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49852),
            .ce(),
            .sr(N__49539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_10_25_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_10_25_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_10_25_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_10_25_2  (
            .in0(N__43129),
            .in1(N__28783),
            .in2(_gnd_net_),
            .in3(N__26611),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49852),
            .ce(),
            .sr(N__49539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_10_25_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_10_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_10_25_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_10_25_3  (
            .in0(N__43137),
            .in1(N__29143),
            .in2(_gnd_net_),
            .in3(N__26608),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49852),
            .ce(),
            .sr(N__49539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_10_25_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_10_25_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_10_25_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_10_25_4  (
            .in0(N__43130),
            .in1(N__29155),
            .in2(_gnd_net_),
            .in3(N__26605),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49852),
            .ce(),
            .sr(N__49539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_10_25_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_10_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_10_25_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_10_25_5  (
            .in0(N__43138),
            .in1(N__29088),
            .in2(_gnd_net_),
            .in3(N__26602),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49852),
            .ce(),
            .sr(N__49539));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_10_25_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_10_25_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_10_25_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_10_25_6  (
            .in0(N__43131),
            .in1(N__29114),
            .in2(_gnd_net_),
            .in3(N__26599),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49852),
            .ce(),
            .sr(N__49539));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_11_4_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_11_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIGC8D_3_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34774),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_11_4_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_11_4_6 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNID56U_7_LC_11_4_6  (
            .in0(N__37983),
            .in1(N__34775),
            .in2(N__33463),
            .in3(N__30121),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNID56UZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_11_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_11_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIIE8D_5_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29614),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_11_5_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_11_5_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_11_5_2 .LUT_INIT=16'b0000101100011011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_11_5_2  (
            .in0(N__37707),
            .in1(N__37499),
            .in2(N__26629),
            .in3(N__37303),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49953),
            .ce(),
            .sr(N__49415));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_11_5_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_11_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILH8D_8_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37091),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_11_6_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_11_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CRY_0_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__29652),
            .in2(N__29656),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_6_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_0_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__29373),
            .in2(N__29356),
            .in3(N__26719),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0_c_THRU_CO ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_6_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_1_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__26716),
            .in2(N__29389),
            .in3(N__26698),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_6_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__26695),
            .in2(N__29224),
            .in3(N__26680),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_6_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__26677),
            .in2(N__26668),
            .in3(N__26656),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_6_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__26653),
            .in2(N__29533),
            .in3(N__26641),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_6_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__29593),
            .in2(N__26638),
            .in3(N__26617),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_6_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__26818),
            .in2(N__29290),
            .in3(N__26797),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_7_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__26794),
            .in2(N__29164),
            .in3(N__26782),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_7_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__26779),
            .in2(N__35146),
            .in3(N__26770),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_7_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__35599),
            .in2(N__29281),
            .in3(N__26767),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_7_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__29503),
            .in2(N__29524),
            .in3(N__26764),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_7_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__27103),
            .in2(N__35230),
            .in3(N__26755),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_7_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__26752),
            .in2(N__29755),
            .in3(N__26734),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_7_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__29497),
            .in2(N__29512),
            .in3(N__26731),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_7_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__26932),
            .in2(N__29173),
            .in3(N__26917),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_8_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__26914),
            .in2(N__29443),
            .in3(N__26896),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_8_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__35317),
            .in2(N__37729),
            .in3(N__26893),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_8_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__33676),
            .in2(N__29665),
            .in3(N__26884),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_8_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__26881),
            .in2(N__35056),
            .in3(N__26860),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_8_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__35608),
            .in2(N__29746),
            .in3(N__26848),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_8_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__29938),
            .in2(N__29947),
            .in3(N__26845),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_8_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__29725),
            .in2(N__33769),
            .in3(N__26842),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_8_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__29803),
            .in2(N__26839),
            .in3(N__27049),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__27394),
            .in2(N__29956),
            .in3(N__27037),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__34120),
            .in2(N__35398),
            .in3(N__27022),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__27079),
            .in2(N__29737),
            .in3(N__27019),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__27073),
            .in2(N__29677),
            .in3(N__27007),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__34039),
            .in2(N__27004),
            .in3(N__26983),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__27092),
            .in2(N__27112),
            .in3(N__26974),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__27094),
            .in2(N__27157),
            .in3(N__26965),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__27093),
            .in2(N__26962),
            .in3(N__26935),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un13_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un13_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_10_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_11_10_0  (
            .in0(N__37460),
            .in1(N__37838),
            .in2(_gnd_net_),
            .in3(N__27205),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI8OI5_29_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27189),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_10_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7NI5_28_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27140),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_11_10_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_11_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVDH5_11_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35273),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_10_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_14_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37837),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_11_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_11_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4KI5_25_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30291),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_11_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_11_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5LI5_26_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29704),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_11_3.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_11_3.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_11_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_11_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27064),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49920),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_11_5 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_11_5  (
            .in0(N__35365),
            .in1(N__29055),
            .in2(_gnd_net_),
            .in3(N__28997),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_400_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_11_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_11_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI2II5_23_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29999),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_12_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_12_2  (
            .in0(N__27385),
            .in1(N__27856),
            .in2(_gnd_net_),
            .in3(N__32850),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_11_12_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27376),
            .in3(N__30257),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49914),
            .ce(),
            .sr(N__49462));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32851),
            .lcout(\current_shift_inst.N_1474_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_12_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_11_12_7  (
            .in0(N__32852),
            .in1(N__27373),
            .in2(_gnd_net_),
            .in3(N__27829),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_13_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_11_13_0  (
            .in0(N__28351),
            .in1(N__27364),
            .in2(_gnd_net_),
            .in3(N__32848),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_13_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_11_13_4  (
            .in0(N__31957),
            .in1(N__27348),
            .in2(N__32668),
            .in3(N__27304),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_14_0 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_11_14_0  (
            .in0(N__27280),
            .in1(N__32445),
            .in2(N__27238),
            .in3(N__31956),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_14_1 .LUT_INIT=16'b1100010111000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_11_14_1  (
            .in0(N__27279),
            .in1(N__27234),
            .in2(N__32025),
            .in3(N__32446),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_11_14_2  (
            .in0(N__27670),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49905),
            .ce(N__27632),
            .sr(N__49478));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_14_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_11_14_3  (
            .in0(N__31952),
            .in1(N__32447),
            .in2(N__27574),
            .in3(N__27601),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_11_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_11_14_4 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_11_14_4  (
            .in0(N__27600),
            .in1(N__27570),
            .in2(N__32588),
            .in3(N__31950),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_14_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_11_14_5  (
            .in0(N__31951),
            .in1(N__27502),
            .in2(_gnd_net_),
            .in3(N__27493),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27532),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_11_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_11_14_7 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_11_14_7  (
            .in0(N__31949),
            .in1(_gnd_net_),
            .in2(N__27496),
            .in3(N__27492),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__27924),
            .in2(N__27460),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_15_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_11_15_1  (
            .in0(N__27991),
            .in1(N__27418),
            .in2(N__27451),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__32318),
            .in2(N__27727),
            .in3(N__27990),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__30772),
            .in2(N__32522),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__32322),
            .in2(N__27718),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__30691),
            .in2(N__32523),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__32326),
            .in2(N__27706),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__27691),
            .in2(N__32524),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__32346),
            .in2(N__27679),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__30946),
            .in2(N__32529),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__32350),
            .in2(N__31378),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__27775),
            .in2(N__32530),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__32354),
            .in2(N__27766),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__30865),
            .in2(N__32531),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__32358),
            .in2(N__31282),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__27757),
            .in2(N__32532),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__32537),
            .in2(N__27751),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__27742),
            .in2(N__32646),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__32541),
            .in2(N__27736),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__31759),
            .in2(N__32647),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__32545),
            .in2(N__27871),
            .in3(N__27844),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__27841),
            .in2(N__32648),
            .in3(N__27820),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__32549),
            .in2(N__31198),
            .in3(N__27817),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__31489),
            .in2(N__32649),
            .in3(N__27814),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__32553),
            .in2(N__31576),
            .in3(N__27811),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__27808),
            .in2(N__32650),
            .in3(N__27802),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__32557),
            .in2(N__27799),
            .in3(N__27790),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__27787),
            .in2(N__32651),
            .in3(N__27778),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__32561),
            .in2(N__28387),
            .in3(N__28372),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__28369),
            .in2(N__32652),
            .in3(N__28363),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__32565),
            .in2(N__28360),
            .in3(N__28342),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_18_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_11_18_7  (
            .in0(N__28339),
            .in1(N__28327),
            .in2(N__32849),
            .in3(N__28318),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_11_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_11_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_11_19_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_11_19_0  (
            .in0(N__47112),
            .in1(N__34518),
            .in2(_gnd_net_),
            .in3(N__42213),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49873),
            .ce(N__49120),
            .sr(N__49511));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_11_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_11_19_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_11_19_2  (
            .in0(N__28220),
            .in1(N__27972),
            .in2(_gnd_net_),
            .in3(N__27943),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__33166),
            .in2(N__27904),
            .in3(N__28719),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_11_20_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(N__27877),
            .in2(N__31726),
            .in3(N__27895),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(N__31747),
            .in2(N__28564),
            .in3(N__28579),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__28540),
            .in2(N__31714),
            .in3(N__28555),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_11_20_4  (
            .in0(_gnd_net_),
            .in1(N__31702),
            .in2(N__28519),
            .in3(N__28534),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(N__31735),
            .in2(N__28492),
            .in3(N__28507),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_20_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_11_20_6  (
            .in0(N__28483),
            .in1(N__28468),
            .in2(N__33175),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_20_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_11_20_7  (
            .in0(N__28462),
            .in1(N__32734),
            .in2(N__28447),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(N__43165),
            .in2(N__28420),
            .in3(N__28438),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_11_21_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(N__43276),
            .in2(N__28396),
            .in3(N__28411),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__43234),
            .in2(N__28681),
            .in3(N__28696),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(N__43195),
            .in2(N__28657),
            .in3(N__28672),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_11_21_4  (
            .in0(_gnd_net_),
            .in1(N__43180),
            .in2(N__28633),
            .in3(N__28648),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_21_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_11_21_5  (
            .in0(N__28624),
            .in1(N__43324),
            .in2(N__28609),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_21_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_11_21_6  (
            .in0(N__28600),
            .in1(N__28585),
            .in2(N__34684),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_21_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_11_21_7  (
            .in0(_gnd_net_),
            .in1(N__42661),
            .in2(N__42739),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_22_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__28891),
            .in2(N__42820),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_22_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_22_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__28858),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_22_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_22_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__28825),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_22_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_22_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_11_22_3  (
            .in0(_gnd_net_),
            .in1(N__28792),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_22_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_22_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_11_22_4  (
            .in0(_gnd_net_),
            .in1(N__28759),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_22_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_22_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__29131),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_22_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__29068),
            .in2(N__29122),
            .in3(N__28750),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28747),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_LC_11_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_11_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_11_23_0 .LUT_INIT=16'b1100010011101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_11_23_0  (
            .in0(N__28920),
            .in1(N__28732),
            .in2(N__28906),
            .in3(N__33086),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(N__49527));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_11_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_11_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1_28_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__28919),
            .in2(_gnd_net_),
            .in3(N__28938),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIM9HS1Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_23_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_23_2 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_11_23_2  (
            .in0(N__33061),
            .in1(N__33084),
            .in2(_gnd_net_),
            .in3(N__28731),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_hc.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_23_3 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_11_23_3  (
            .in0(N__43042),
            .in1(N__28939),
            .in2(N__28723),
            .in3(N__28718),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(N__49527));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_11_23_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_11_23_4 .LUT_INIT=16'b1101110011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI1LP11_28_LC_11_23_4  (
            .in0(N__29089),
            .in1(N__29115),
            .in2(N__28951),
            .in3(N__33085),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_23_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28930),
            .in3(N__28918),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_11_23_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_11_23_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_11_23_6 .LUT_INIT=16'b1101110100001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_11_23_6  (
            .in0(N__28921),
            .in1(N__33087),
            .in2(N__28905),
            .in3(N__44624),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49856),
            .ce(),
            .sr(N__49527));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_11_24_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_11_24_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_11_24_1  (
            .in0(N__43345),
            .in1(N__42866),
            .in2(N__42846),
            .in3(N__42898),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_24_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_24_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_11_24_2  (
            .in0(_gnd_net_),
            .in1(N__28881),
            .in2(_gnd_net_),
            .in3(N__28869),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_11_24_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_11_24_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_11_24_3  (
            .in0(N__28848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28836),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_11_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_11_24_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_11_24_4  (
            .in0(_gnd_net_),
            .in1(N__28815),
            .in2(_gnd_net_),
            .in3(N__28803),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_24_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_24_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_11_24_5  (
            .in0(_gnd_net_),
            .in1(N__28782),
            .in2(_gnd_net_),
            .in3(N__28770),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_24_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_24_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_24_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(N__29154),
            .in2(_gnd_net_),
            .in3(N__29142),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_df28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_24_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_24_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_11_24_7  (
            .in0(_gnd_net_),
            .in1(N__29113),
            .in2(_gnd_net_),
            .in3(N__29087),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_25_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_25_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_25_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_11_25_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29048),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29020),
            .ce(),
            .sr(N__49536));
    defparam \delay_measurement_inst.start_timer_tr_LC_11_26_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_11_26_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_11_26_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_11_26_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29047),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29019),
            .ce(),
            .sr(N__49540));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_3_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_3_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__35383),
            .in2(_gnd_net_),
            .in3(N__29008),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_399_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_4_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIV7J_7_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30120),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_4_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIU6J_6_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30146),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_4_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIS4J_4_LC_12_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29912),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_4_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIT5J_5_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29882),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_5_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI5R3U_5_LC_12_5_1  (
            .in0(N__37878),
            .in1(N__29430),
            .in2(N__29887),
            .in3(N__33184),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI5R3UZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_12_5_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_12_5_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1M2U_4_LC_12_5_2  (
            .in0(N__29377),
            .in1(N__37877),
            .in2(N__29917),
            .in3(N__33199),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI1M2UZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_12_5_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_12_5_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI7T941_10_LC_12_5_3  (
            .in0(N__37882),
            .in1(N__29339),
            .in2(N__33415),
            .in3(N__30057),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI7T941Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_12_5_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_12_5_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIQ6T01_13_LC_12_5_4  (
            .in0(N__38096),
            .in1(N__37883),
            .in2(N__33754),
            .in3(N__33376),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIQ6T01Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_12_5_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_12_5_5 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI905U_6_LC_12_5_5  (
            .in0(N__29266),
            .in1(N__30147),
            .in2(N__37942),
            .in3(N__33478),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNI905UZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_5_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_5_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI09J_8_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30086),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_5_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI9FJ3_10_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30056),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_12_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_12_6_0 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4I_LC_12_6_0  (
            .in0(N__33546),
            .in1(N__29214),
            .in2(N__33529),
            .in3(N__37974),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_RNIJA4IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_12_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_12_6_1 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIISQ01_11_LC_12_6_1  (
            .in0(N__37972),
            .in1(N__33951),
            .in2(N__33394),
            .in3(N__30033),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIISQ01Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_12_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_12_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIDJJ3_0_14_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37969),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_12_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_12_6_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNILF8U_9_LC_12_6_3  (
            .in0(N__37971),
            .in1(N__29623),
            .in2(N__33433),
            .in3(N__35020),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNILF8UZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_12_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_12_6_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIHA7U_8_LC_12_6_4  (
            .in0(N__29583),
            .in1(N__37970),
            .in2(N__30091),
            .in3(N__33442),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIHA7UZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIAGJ3_11_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30032),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_12_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_12_6_6 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVH_LC_12_6_6  (
            .in0(N__35041),
            .in1(N__33867),
            .in2(N__33583),
            .in3(N__37973),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_c_RNIBUVHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_12_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_12_7_0 .LUT_INIT=16'b0111110101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73I_LC_12_7_0  (
            .in0(N__37871),
            .in1(N__33556),
            .in2(N__35494),
            .in3(N__38155),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_RNIH73IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_12_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_12_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUCH5_10_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33840),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1GH5_13_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38154),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_12_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_12_7_3 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5I_LC_12_7_3  (
            .in0(N__34987),
            .in1(N__29491),
            .in2(N__33514),
            .in3(N__37872),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_RNILD5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_12_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_12_7_4 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96J_LC_12_7_4  (
            .in0(N__29856),
            .in1(N__35515),
            .in2(N__37941),
            .in3(N__33622),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_RNIH96JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_c_inv_LC_12_7_5  (
            .in0(N__33547),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37867),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_12_7_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_12_7_6 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42I_LC_12_7_6  (
            .in0(N__29789),
            .in1(N__34144),
            .in2(N__37940),
            .in3(N__33565),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_RNIF42IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_12_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_12_7_7 .LUT_INIT=16'b0101101011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82J_LC_12_7_7  (
            .in0(N__35215),
            .in1(N__35650),
            .in2(N__33664),
            .in3(N__37873),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_RNIK82JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_12_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_12_8_0 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9J_LC_12_8_0  (
            .in0(N__30311),
            .in1(N__34177),
            .in2(N__37944),
            .in3(N__33601),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_RNINI9JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_c_inv_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(N__33643),
            .in2(_gnd_net_),
            .in3(N__37884),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_12_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_12_8_2 .LUT_INIT=16'b0111110101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65J_LC_12_8_2  (
            .in0(N__37888),
            .in1(N__33631),
            .in2(N__29728),
            .in3(N__33802),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_RNIF65JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_12_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_12_8_3 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJ_LC_12_8_3  (
            .in0(N__29719),
            .in1(N__37892),
            .in2(N__35587),
            .in3(N__33592),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_RNIPLAJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_12_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_12_8_4 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20J_LC_12_8_4  (
            .in0(N__33716),
            .in1(N__35341),
            .in2(N__37943),
            .in3(N__33499),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_RNIG20JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_12_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_12_8_5 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7J_LC_12_8_5  (
            .in0(N__34109),
            .in1(N__30004),
            .in2(N__37945),
            .in3(N__33613),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_RNIJC7JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_12_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_12_8_6 .LUT_INIT=16'b0111011110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34J_LC_12_8_6  (
            .in0(N__35308),
            .in1(N__37893),
            .in2(N__34011),
            .in3(N__33652),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_RNID34JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVEI5_20_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34002),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_9_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__29932),
            .in2(_gnd_net_),
            .in3(N__30235),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_9_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_9_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_12_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__30220),
            .in2(_gnd_net_),
            .in3(N__29926),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__49925),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_9_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_12_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__30208),
            .in2(_gnd_net_),
            .in3(N__29923),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__49925),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_9_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_12_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__30196),
            .in2(_gnd_net_),
            .in3(N__29920),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__49925),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_9_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_9_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_12_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__30184),
            .in2(_gnd_net_),
            .in3(N__29890),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__49925),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_9_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_9_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_12_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(N__30172),
            .in2(_gnd_net_),
            .in3(N__29860),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__49925),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_9_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_9_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_12_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__30160),
            .in2(_gnd_net_),
            .in3(N__30124),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__49925),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_9_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_9_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_12_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(N__30451),
            .in2(_gnd_net_),
            .in3(N__30094),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__49925),
            .ce(),
            .sr(N__49431));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_10_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_10_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_12_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__30439),
            .in2(_gnd_net_),
            .in3(N__30064),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__49918),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_10_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_12_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__30427),
            .in2(_gnd_net_),
            .in3(N__30061),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__49918),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_10_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_12_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__30409),
            .in2(_gnd_net_),
            .in3(N__30037),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__49918),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_10_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_12_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__30385),
            .in2(_gnd_net_),
            .in3(N__30013),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__49918),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_10_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_12_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__30364),
            .in2(_gnd_net_),
            .in3(N__30010),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__49918),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_12_10_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_12_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(N__30337),
            .in2(_gnd_net_),
            .in3(N__30007),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__49918),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_12_10_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_12_10_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(N__30349),
            .in2(_gnd_net_),
            .in3(N__30328),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_12_10_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_12_10_7 .LUT_INIT=16'b0010111100101110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_12_10_7  (
            .in0(N__37475),
            .in1(N__37681),
            .in2(N__30325),
            .in3(N__37316),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49918),
            .ce(),
            .sr(N__49438));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__30268),
            .in2(N__30261),
            .in3(N__30262),
            .lcout(\current_shift_inst.control_input_18 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__30226),
            .in2(_gnd_net_),
            .in3(N__30211),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__31672),
            .in2(_gnd_net_),
            .in3(N__30199),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__33022),
            .in2(_gnd_net_),
            .in3(N__30187),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__32992),
            .in2(_gnd_net_),
            .in3(N__30175),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__32962),
            .in2(_gnd_net_),
            .in3(N__30163),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__32935),
            .in2(_gnd_net_),
            .in3(N__30151),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__32905),
            .in2(_gnd_net_),
            .in3(N__30442),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__32749),
            .in2(_gnd_net_),
            .in3(N__30430),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__31465),
            .in2(_gnd_net_),
            .in3(N__30418),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__30415),
            .in2(_gnd_net_),
            .in3(N__30400),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__30397),
            .in2(_gnd_net_),
            .in3(N__30376),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__30373),
            .in2(_gnd_net_),
            .in3(N__30355),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__32857),
            .in2(_gnd_net_),
            .in3(N__30352),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(\current_shift_inst.control_input_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30340),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_0_LC_12_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_12_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_12_13_0 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst2.state_0_LC_12_13_0  (
            .in0(N__30669),
            .in1(N__35844),
            .in2(N__30685),
            .in3(N__35873),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49904),
            .ce(),
            .sr(N__49463));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_12_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_12_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__30668),
            .in2(_gnd_net_),
            .in3(N__30681),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_12_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_12_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_12_13_2 .LUT_INIT=16'b1100010011110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_12_13_2  (
            .in0(N__35794),
            .in1(N__36229),
            .in2(N__30673),
            .in3(N__36141),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49904),
            .ce(),
            .sr(N__49463));
    defparam \phase_controller_inst2.state_1_LC_12_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_12_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_12_13_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst2.state_1_LC_12_13_3  (
            .in0(N__35845),
            .in1(N__35872),
            .in2(_gnd_net_),
            .in3(N__41278),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49904),
            .ce(),
            .sr(N__49463));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_13_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_13_5  (
            .in0(N__36140),
            .in1(N__36106),
            .in2(N__36078),
            .in3(N__36739),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49904),
            .ce(),
            .sr(N__49463));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_12_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_12_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_12_14_0 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_12_14_0  (
            .in0(N__35740),
            .in1(N__38793),
            .in2(N__38860),
            .in3(N__40696),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49899),
            .ce(N__50321),
            .sr(N__49470));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_12_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_12_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_12_14_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_12_14_1  (
            .in0(N__38792),
            .in1(N__41803),
            .in2(_gnd_net_),
            .in3(N__35719),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49899),
            .ce(N__50321),
            .sr(N__49470));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_12_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_12_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_12_14_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_12_14_2  (
            .in0(N__41804),
            .in1(N__35683),
            .in2(_gnd_net_),
            .in3(N__38794),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49899),
            .ce(N__50321),
            .sr(N__49470));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_12_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_12_14_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_12_14_6  (
            .in0(N__30658),
            .in1(N__30531),
            .in2(_gnd_net_),
            .in3(N__30486),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_12_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_12_15_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_12_15_0  (
            .in0(N__32451),
            .in1(N__31964),
            .in2(N__31189),
            .in3(N__31138),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_15_2 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_12_15_2  (
            .in0(N__32453),
            .in1(N__31961),
            .in2(N__31095),
            .in3(N__31058),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_12_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_12_15_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_12_15_3  (
            .in0(N__31960),
            .in1(N__32457),
            .in2(N__31015),
            .in3(N__30970),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_15_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_12_15_4  (
            .in0(N__32452),
            .in1(N__31962),
            .in2(N__30940),
            .in3(N__30892),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_12_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_12_15_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_12_15_5  (
            .in0(N__31963),
            .in1(N__32454),
            .in2(N__31804),
            .in3(N__31830),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_12_15_6  (
            .in0(N__32455),
            .in1(N__31958),
            .in2(N__30849),
            .in3(N__30799),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_12_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_12_15_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_12_15_7  (
            .in0(N__31959),
            .in1(N__32456),
            .in2(N__30766),
            .in3(N__30718),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36180),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49887),
            .ce(),
            .sr(N__49485));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_16_5 .LUT_INIT=16'b1101110000001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_12_16_5  (
            .in0(N__50058),
            .in1(N__34649),
            .in2(N__50037),
            .in3(N__50107),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49887),
            .ce(),
            .sr(N__49485));
    defparam \phase_controller_inst1.state_4_LC_12_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_12_16_6 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_12_16_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_12_16_6  (
            .in0(N__33140),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44532),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49887),
            .ce(),
            .sr(N__49485));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_12_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_12_17_0 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_12_17_0  (
            .in0(N__32137),
            .in1(N__31657),
            .in2(N__31608),
            .in3(N__32594),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_17_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_12_17_1  (
            .in0(N__32593),
            .in1(N__32136),
            .in2(N__31563),
            .in3(N__31516),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_12_17_2  (
            .in0(N__31483),
            .in1(N__31477),
            .in2(_gnd_net_),
            .in3(N__32828),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_17_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_12_17_3  (
            .in0(N__32595),
            .in1(N__32132),
            .in2(N__31456),
            .in3(N__31419),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_12_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_12_17_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_12_17_4  (
            .in0(N__32133),
            .in1(N__32596),
            .in2(N__31368),
            .in3(N__31312),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_17_5 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_12_17_5  (
            .in0(N__32592),
            .in1(N__32135),
            .in2(N__31273),
            .in3(N__31239),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_12_17_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_12_17_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9AJ01_27_LC_12_17_6  (
            .in0(N__39516),
            .in1(N__42547),
            .in2(N__39493),
            .in3(N__42525),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_17_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_12_17_7  (
            .in0(N__32597),
            .in1(N__32134),
            .in2(N__31837),
            .in3(N__31803),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_12_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_12_18_0 .LUT_INIT=16'b1110111011111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFKEE1_3_LC_12_18_0  (
            .in0(N__46015),
            .in1(N__39241),
            .in2(N__34609),
            .in3(N__45547),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_12_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_12_18_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRB3CP1_3_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31753),
            .in3(N__45370),
            .lcout(elapsed_time_ns_1_RNIRB3CP1_0_3),
            .ltout(elapsed_time_ns_1_RNIRB3CP1_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_12_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_12_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_12_18_2 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_12_18_2  (
            .in0(N__42280),
            .in1(N__42201),
            .in2(N__31750),
            .in3(N__34483),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(N__43150),
            .sr(N__49500));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_12_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_12_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_12_18_3 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_12_18_3  (
            .in0(N__47088),
            .in1(N__45964),
            .in2(N__42215),
            .in3(N__42283),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(N__43150),
            .sr(N__49500));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_12_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_12_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_12_18_4 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_12_18_4  (
            .in0(N__42279),
            .in1(N__47085),
            .in2(N__34702),
            .in3(N__42200),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(N__43150),
            .sr(N__49500));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_12_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_12_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_12_18_5 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_12_18_5  (
            .in0(N__47086),
            .in1(N__42282),
            .in2(N__42214),
            .in3(N__39303),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(N__43150),
            .sr(N__49500));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_12_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_12_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_12_18_6 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_12_18_6  (
            .in0(N__42281),
            .in1(N__47087),
            .in2(N__42313),
            .in3(N__42202),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49872),
            .ce(N__43150),
            .sr(N__49500));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_19_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_19_0  (
            .in0(N__31693),
            .in1(N__31681),
            .in2(_gnd_net_),
            .in3(N__32821),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_19_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_19_1  (
            .in0(N__32823),
            .in1(N__33043),
            .in2(_gnd_net_),
            .in3(N__33031),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_19_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_19_2  (
            .in0(N__33010),
            .in1(N__32998),
            .in2(_gnd_net_),
            .in3(N__32824),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_19_3 .LUT_INIT=16'b0010011100100111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_19_3  (
            .in0(N__32826),
            .in1(N__32983),
            .in2(N__32977),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_19_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_19_4  (
            .in0(N__32953),
            .in1(N__32947),
            .in2(_gnd_net_),
            .in3(N__32822),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_19_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_19_5  (
            .in0(N__32825),
            .in1(N__32923),
            .in2(_gnd_net_),
            .in3(N__32917),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_19_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32893),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_19_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_19_7  (
            .in0(N__32827),
            .in1(N__32767),
            .in2(_gnd_net_),
            .in3(N__32755),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_12_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_12_20_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_12_20_0  (
            .in0(N__47098),
            .in1(N__42204),
            .in2(_gnd_net_),
            .in3(N__34519),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(N__43144),
            .sr(N__49512));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_12_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_12_20_4 .LUT_INIT=16'b0100000001000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_12_20_4  (
            .in0(N__47097),
            .in1(N__42203),
            .in2(N__38323),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(N__43144),
            .sr(N__49512));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_12_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_12_20_6 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_12_20_6  (
            .in0(N__34534),
            .in1(N__42284),
            .in2(N__34720),
            .in3(N__34735),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49862),
            .ce(N__43144),
            .sr(N__49512));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_21_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(N__38246),
            .in2(_gnd_net_),
            .in3(N__38295),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_12_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_12_21_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a2_1_LC_12_21_3  (
            .in0(N__33149),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44541),
            .lcout(state_ns_i_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_12_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_12_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_12_22_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_12_22_2  (
            .in0(N__33066),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(N__49522));
    defparam \phase_controller_inst1.state_1_LC_12_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_12_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_12_22_5 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \phase_controller_inst1.state_1_LC_12_22_5  (
            .in0(N__33367),
            .in1(N__44601),
            .in2(_gnd_net_),
            .in3(N__46643),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(N__49522));
    defparam \phase_controller_inst1.start_timer_hc_LC_12_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_12_22_6 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_12_22_6  (
            .in0(N__44542),
            .in1(N__33366),
            .in2(N__33067),
            .in3(N__33094),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49854),
            .ce(),
            .sr(N__49522));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_23_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__33088),
            .in2(_gnd_net_),
            .in3(N__33062),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_23_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_12_23_1  (
            .in0(N__34659),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34918),
            .lcout(\phase_controller_inst1.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_12_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_12_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(N__46598),
            .in2(_gnd_net_),
            .in3(N__44618),
            .lcout(\phase_controller_inst1.N_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_24_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_12_24_2  (
            .in0(N__34957),
            .in1(N__34877),
            .in2(_gnd_net_),
            .in3(N__34850),
            .lcout(\current_shift_inst.timer_s1.N_167_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_4_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_0_c_inv_LC_13_4_0  (
            .in0(_gnd_net_),
            .in1(N__33295),
            .in2(_gnd_net_),
            .in3(N__33316),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_0 ),
            .ltout(),
            .carryin(bfn_13_4_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_4_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_1_c_inv_LC_13_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33268),
            .in3(N__33289),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_4_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_2_c_inv_LC_13_4_2  (
            .in0(_gnd_net_),
            .in1(N__33238),
            .in2(_gnd_net_),
            .in3(N__33259),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_4_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_4_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_inv_LC_13_4_3  (
            .in0(_gnd_net_),
            .in1(N__33211),
            .in2(_gnd_net_),
            .in3(N__33232),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_4_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_4_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_3_c_RNIBKJC_LC_13_4_4  (
            .in0(_gnd_net_),
            .in1(N__33205),
            .in2(_gnd_net_),
            .in3(N__33193),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_4_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_4_c_RNIDNKC_LC_13_4_5  (
            .in0(_gnd_net_),
            .in1(N__33190),
            .in2(_gnd_net_),
            .in3(N__33178),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_4_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_5_c_RNIFQLC_LC_13_4_6  (
            .in0(_gnd_net_),
            .in1(N__33484),
            .in2(_gnd_net_),
            .in3(N__33472),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_4_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_4_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_6_c_RNIHTMC_LC_13_4_7  (
            .in0(_gnd_net_),
            .in1(N__33469),
            .in2(_gnd_net_),
            .in3(N__33451),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_5_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_7_c_RNIJ0OC_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(N__33448),
            .in2(_gnd_net_),
            .in3(N__33436),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_8 ),
            .ltout(),
            .carryin(bfn_13_5_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_5_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_8_c_RNIL3PC_LC_13_5_1  (
            .in0(_gnd_net_),
            .in1(N__34993),
            .in2(_gnd_net_),
            .in3(N__33424),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_5_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_9_c_RNIUAQF_LC_13_5_2  (
            .in0(_gnd_net_),
            .in1(N__33421),
            .in2(_gnd_net_),
            .in3(N__33403),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_5_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_10_c_RNI78BC_LC_13_5_3  (
            .in0(_gnd_net_),
            .in1(N__33400),
            .in2(_gnd_net_),
            .in3(N__33382),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_13_5_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_13_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_11_c_RNI9BCC_LC_13_5_4  (
            .in0(_gnd_net_),
            .in1(N__34753),
            .in2(_gnd_net_),
            .in3(N__33379),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_13_5_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_13_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_12_c_RNIBEDC_LC_13_5_5  (
            .in0(_gnd_net_),
            .in1(N__33727),
            .in2(_gnd_net_),
            .in3(N__33370),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_5_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_LUT4_0_LC_13_5_6  (
            .in0(_gnd_net_),
            .in1(N__35036),
            .in2(_gnd_net_),
            .in3(N__33571),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_5_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_LUT4_0_LC_13_5_7  (
            .in0(_gnd_net_),
            .in1(N__34746),
            .in2(_gnd_net_),
            .in3(N__33568),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_6_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_LUT4_0_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__34140),
            .in2(_gnd_net_),
            .in3(N__33559),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_6_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_LUT4_0_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__35486),
            .in2(_gnd_net_),
            .in3(N__33550),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_6_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_LUT4_0_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__33545),
            .in2(_gnd_net_),
            .in3(N__33517),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_6_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_LUT4_0_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__34979),
            .in2(_gnd_net_),
            .in3(N__33505),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_6_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_LUT4_0_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__38057),
            .in2(_gnd_net_),
            .in3(N__33502),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_6_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_LUT4_0_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__35340),
            .in2(_gnd_net_),
            .in3(N__33490),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_6_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_LUT4_0_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__35078),
            .in2(_gnd_net_),
            .in3(N__33487),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_6_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_LUT4_0_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__35207),
            .in2(_gnd_net_),
            .in3(N__33655),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_7_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_LUT4_0_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35307),
            .in3(N__33646),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_THRU_CO ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_7_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_LUT4_0_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__33642),
            .in2(_gnd_net_),
            .in3(N__33625),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_7_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_LUT4_0_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__35510),
            .in2(_gnd_net_),
            .in3(N__33616),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_7_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_LUT4_0_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__34111),
            .in2(_gnd_net_),
            .in3(N__33607),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_7_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_LUT4_0_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__35469),
            .in2(_gnd_net_),
            .in3(N__33604),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_7_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_LUT4_0_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__34173),
            .in2(_gnd_net_),
            .in3(N__33595),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_7_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_LUT4_0_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(N__35579),
            .in2(_gnd_net_),
            .in3(N__33586),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un7_integrator1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_13_7_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_13_7_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74K_LC_13_7_7  (
            .in0(N__34086),
            .in1(N__37946),
            .in2(_gnd_net_),
            .in3(N__34042),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_RNII74KZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_13_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_13_8_2 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_13_8_2  (
            .in0(N__37287),
            .in1(N__37495),
            .in2(N__34027),
            .in3(N__37612),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49420));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_13_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_13_8_4 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_13_8_4  (
            .in0(N__37288),
            .in1(N__37496),
            .in2(N__33979),
            .in3(N__37613),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49420));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_13_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_13_8_5 .LUT_INIT=16'b0000000111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_13_8_5  (
            .in0(N__37493),
            .in1(N__37290),
            .in2(N__37668),
            .in3(N__33967),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49420));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_13_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_13_8_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_13_8_6 .LUT_INIT=16'b0000111111001110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_13_8_6  (
            .in0(N__37286),
            .in1(N__37494),
            .in2(N__33895),
            .in3(N__37614),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49420));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_13_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_13_8_7 .LUT_INIT=16'b0000101011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_13_8_7  (
            .in0(N__37492),
            .in1(N__37289),
            .in2(N__37667),
            .in3(N__33883),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49938),
            .ce(),
            .sr(N__49420));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_13_9_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_13_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI0GI5_21_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33792),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNICIJ3_13_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33743),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_13_9_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_13_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5KH5_17_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33717),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_16_c_inv_LC_13_9_4  (
            .in0(N__34139),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37791),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_13_9_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_13_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI3JI5_24_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35442),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_13_9_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_13_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_inv_LC_13_9_7  (
            .in0(N__37792),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34110),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_13_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_13_10_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_13_10_1  (
            .in0(N__41634),
            .in1(N__38427),
            .in2(N__38500),
            .in3(N__41808),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49926),
            .ce(N__36763),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_13_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_13_10_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_13_10_2  (
            .in0(N__41807),
            .in1(N__38522),
            .in2(N__38431),
            .in3(N__41637),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49926),
            .ce(N__36763),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_13_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_13_10_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_13_10_3  (
            .in0(N__41633),
            .in1(N__38426),
            .in2(N__38572),
            .in3(N__41805),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49926),
            .ce(N__36763),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_13_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_13_10_5 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_13_10_5  (
            .in0(N__41635),
            .in1(N__41809),
            .in2(N__41449),
            .in3(N__38428),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49926),
            .ce(N__36763),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_13_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_13_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_13_10_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_13_10_6  (
            .in0(N__41806),
            .in1(N__38547),
            .in2(N__38430),
            .in3(N__41636),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49926),
            .ce(N__36763),
            .sr(N__49432));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_11_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__36817),
            .in2(_gnd_net_),
            .in3(N__36838),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__37050),
            .in2(_gnd_net_),
            .in3(N__36796),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_13_11_2 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_13_11_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_13_11_2  (
            .in0(N__49583),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_13_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_13_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_29_c_inv_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__34172),
            .in2(_gnd_net_),
            .in3(N__37833),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_13_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_13_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_13_12_0 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_13_12_0  (
            .in0(N__38769),
            .in1(N__41781),
            .in2(N__40642),
            .in3(N__38851),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49915),
            .ce(N__36761),
            .sr(N__49449));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_13_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_13_12_1 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_13_12_1  (
            .in0(N__35733),
            .in1(N__38844),
            .in2(N__38791),
            .in3(N__40692),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49915),
            .ce(N__36761),
            .sr(N__49449));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_13_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_13_12_2 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_13_12_2  (
            .in0(N__38768),
            .in1(N__41779),
            .in2(N__41104),
            .in3(N__38850),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49915),
            .ce(N__36761),
            .sr(N__49449));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_13_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_13_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_13_12_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_13_12_4  (
            .in0(N__35715),
            .in1(N__38776),
            .in2(_gnd_net_),
            .in3(N__41777),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49915),
            .ce(N__36761),
            .sr(N__49449));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_13_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_13_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_13_12_5 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_13_12_5  (
            .in0(N__41780),
            .in1(N__38845),
            .in2(N__41143),
            .in3(N__38770),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49915),
            .ce(N__36761),
            .sr(N__49449));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_13_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_13_12_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_13_12_7  (
            .in0(N__41778),
            .in1(N__35676),
            .in2(_gnd_net_),
            .in3(N__38771),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49915),
            .ce(N__36761),
            .sr(N__49449));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__35752),
            .in2(N__34153),
            .in3(N__36074),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_13_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_13_13_1  (
            .in0(N__36049),
            .in1(N__35746),
            .in2(N__34309),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__34300),
            .in2(N__34294),
            .in3(N__36022),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__34282),
            .in2(N__34276),
            .in3(N__36004),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(N__34267),
            .in2(N__34261),
            .in3(N__35986),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__34249),
            .in2(N__34243),
            .in3(N__36391),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_13_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_13_13_6  (
            .in0(N__36370),
            .in1(N__34225),
            .in2(N__34234),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(N__34210),
            .in2(N__34219),
            .in3(N__36352),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_14_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_13_14_0  (
            .in0(N__36334),
            .in1(N__34204),
            .in2(N__35557),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_13_14_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__34402),
            .in2(N__34414),
            .in3(N__36316),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__34396),
            .in2(N__34387),
            .in3(N__36298),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__34375),
            .in2(N__34366),
            .in3(N__36274),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__34357),
            .in2(N__34348),
            .in3(N__36256),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_13_14_5  (
            .in0(N__36556),
            .in1(N__34336),
            .in2(N__34327),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(N__35542),
            .in2(N__34318),
            .in3(N__36538),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(N__35890),
            .in2(N__35530),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__35941),
            .in2(N__35968),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__36985),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__36943),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__36904),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__36865),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(N__34438),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__34429),
            .in2(N__37057),
            .in3(N__34420),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34417),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_13_16_5  (
            .in0(N__42267),
            .in1(N__34608),
            .in2(N__42220),
            .in3(N__34482),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49894),
            .ce(N__49122),
            .sr(N__49479));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_13_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_13_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHUIH1_10_LC_13_17_0  (
            .in0(N__39340),
            .in1(N__39357),
            .in2(N__45631),
            .in3(N__39372),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_13_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_13_17_1 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPKKEE1_8_LC_13_17_1  (
            .in0(N__39358),
            .in1(N__45560),
            .in2(N__45936),
            .in3(N__34506),
            .lcout(elapsed_time_ns_1_RNIPKKEE1_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_13_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_13_17_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIOJKEE1_7_LC_13_17_2  (
            .in0(N__45929),
            .in1(N__39373),
            .in2(N__45562),
            .in3(N__38312),
            .lcout(elapsed_time_ns_1_RNIOJKEE1_0_7),
            .ltout(elapsed_time_ns_1_RNIOJKEE1_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_13_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_13_17_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_0_2_LC_13_17_3  (
            .in0(N__45959),
            .in1(N__34505),
            .in2(N__34492),
            .in3(N__45786),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_13_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_13_17_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_6_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__46746),
            .in2(N__34489),
            .in3(N__45705),
            .lcout(\phase_controller_inst1.stoper_hc.N_330 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_13_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_13_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_13_17_5 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_13_17_5  (
            .in0(N__45960),
            .in1(N__47084),
            .in2(N__34486),
            .in3(N__42212),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49888),
            .ce(N__49109),
            .sr(N__49486));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_13_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_13_17_7 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_3_LC_13_17_7  (
            .in0(N__46747),
            .in1(N__47083),
            .in2(N__34459),
            .in3(N__34471),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_13_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_13_18_0 .LUT_INIT=16'b0011101100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_0_2_LC_13_18_0  (
            .in0(N__34455),
            .in1(N__34572),
            .in2(N__34607),
            .in3(N__34470),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_13_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_13_18_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJEKEE1_2_LC_13_18_1  (
            .in0(N__34552),
            .in1(N__45937),
            .in2(N__34576),
            .in3(N__45548),
            .lcout(elapsed_time_ns_1_RNIJEKEE1_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_13_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_13_18_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_2_LC_13_18_2  (
            .in0(N__45588),
            .in1(N__46874),
            .in2(N__45730),
            .in3(N__37021),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2 ),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_13_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_13_18_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_a5_1_LC_13_18_3  (
            .in0(N__34561),
            .in1(N__34454),
            .in2(N__34441),
            .in3(N__46800),
            .lcout(\phase_controller_inst1.stoper_hc.N_310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_13_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_13_18_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_o2_1_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__34597),
            .in2(_gnd_net_),
            .in3(N__34571),
            .lcout(\phase_controller_inst1.stoper_hc.N_286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_13_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_13_18_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__46048),
            .in2(_gnd_net_),
            .in3(N__42331),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_13_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_13_18_6 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI63452_2_LC_13_18_6  (
            .in0(N__39223),
            .in1(N__39240),
            .in2(N__34555),
            .in3(N__34551),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_13_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_13_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_13_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39759),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49881),
            .ce(N__39447),
            .sr(N__49492));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_13_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_13_19_0 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0_6_LC_13_19_0  (
            .in0(N__46886),
            .in1(N__45589),
            .in2(_gnd_net_),
            .in3(N__45787),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_13_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_13_19_1 .LUT_INIT=16'b0011001100010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_a2_0_6_LC_13_19_1  (
            .in0(N__45731),
            .in1(N__46812),
            .in2(N__34543),
            .in3(N__45668),
            .lcout(\phase_controller_inst1.stoper_hc.N_328 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_13_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_13_19_2 .LUT_INIT=16'b1100110011111100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_0_0_1_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__47078),
            .in2(N__34540),
            .in3(N__34533),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_0_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_13_19_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_13_19_3 .LUT_INIT=16'b1111001011111110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII3N721_1_LC_13_19_3  (
            .in0(N__34532),
            .in1(N__45561),
            .in2(N__45379),
            .in3(N__39463),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_13_19_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_13_19_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP93CP1_1_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34537),
            .in3(N__46024),
            .lcout(elapsed_time_ns_1_RNIP93CP1_0_1),
            .ltout(elapsed_time_ns_1_RNIP93CP1_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_13_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_13_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_13_19_5 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_13_19_5  (
            .in0(N__42271),
            .in1(N__34734),
            .in2(N__34723),
            .in3(N__34719),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49874),
            .ce(N__49110),
            .sr(N__49501));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_13_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_13_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_13_19_6 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_13_19_6  (
            .in0(N__34701),
            .in1(N__42193),
            .in2(N__42285),
            .in3(N__47079),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49874),
            .ce(N__49110),
            .sr(N__49501));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_13_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_13_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_13_19_7 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_13_19_7  (
            .in0(N__42192),
            .in1(N__42272),
            .in2(N__47105),
            .in3(N__39307),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49874),
            .ce(N__49110),
            .sr(N__49501));
    defparam \phase_controller_inst2.state_3_LC_13_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_13_20_7 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst2.state_3_LC_13_20_7  (
            .in0(N__41246),
            .in1(N__34672),
            .in2(N__41227),
            .in3(N__35818),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49869),
            .ce(),
            .sr(N__49507));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_13_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_13_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_13_21_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_13_21_5  (
            .in0(N__47111),
            .in1(N__46801),
            .in2(N__45736),
            .in3(N__45672),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49864),
            .ce(N__43143),
            .sr(N__49513));
    defparam \phase_controller_inst1.state_3_LC_13_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_13_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_13_22_6 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst1.state_3_LC_13_22_6  (
            .in0(N__38257),
            .in1(N__34671),
            .in2(N__38296),
            .in3(N__44490),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49859),
            .ce(),
            .sr(N__49517));
    defparam \phase_controller_inst1.state_0_LC_13_23_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_13_23_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_13_23_5 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst1.state_0_LC_13_23_5  (
            .in0(N__44602),
            .in1(N__34660),
            .in2(N__46656),
            .in3(N__34920),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49857),
            .ce(),
            .sr(N__49523));
    defparam \phase_controller_inst1.T45_LC_13_23_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.T45_LC_13_23_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T45_LC_13_23_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst1.T45_LC_13_23_7  (
            .in0(N__38254),
            .in1(N__34620),
            .in2(_gnd_net_),
            .in3(N__34919),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49857),
            .ce(),
            .sr(N__49523));
    defparam \current_shift_inst.stop_timer_s1_LC_13_24_0 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_13_24_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_13_24_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_13_24_0  (
            .in0(N__38259),
            .in1(N__34935),
            .in2(N__34963),
            .in3(N__34851),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49853),
            .ce(),
            .sr(N__49525));
    defparam \current_shift_inst.timer_s1.running_LC_13_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_24_1 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_24_1  (
            .in0(N__34852),
            .in1(N__34962),
            .in2(_gnd_net_),
            .in3(N__34878),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49853),
            .ce(),
            .sr(N__49525));
    defparam \current_shift_inst.start_timer_s1_LC_13_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_13_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_13_24_3 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_13_24_3  (
            .in0(N__34934),
            .in1(N__34961),
            .in2(_gnd_net_),
            .in3(N__38258),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49853),
            .ce(),
            .sr(N__49525));
    defparam \phase_controller_inst1.S1_LC_13_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_24_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_13_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38260),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49853),
            .ce(),
            .sr(N__49525));
    defparam \phase_controller_inst1.T23_LC_13_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.T23_LC_13_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T23_LC_13_24_7 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst1.T23_LC_13_24_7  (
            .in0(N__34890),
            .in1(N__46664),
            .in2(_gnd_net_),
            .in3(N__34921),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49853),
            .ce(),
            .sr(N__49525));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_25_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_25_6  (
            .in0(_gnd_net_),
            .in1(N__34873),
            .in2(_gnd_net_),
            .in3(N__34849),
            .lcout(\current_shift_inst.timer_s1.N_166_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S2_LC_13_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_26_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46663),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49850),
            .ce(),
            .sr(N__49532));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_14_4_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_14_4_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_14_4_6 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_14_4_6  (
            .in0(N__37666),
            .in1(N__37323),
            .in2(_gnd_net_),
            .in3(N__34813),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49964),
            .ce(),
            .sr(N__49405));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_5_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIBHJ3_12_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35190),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_14_5_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_14_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_15_c_inv_LC_14_5_1  (
            .in0(N__34747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37976),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_14_5_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_14_5_2 .LUT_INIT=16'b0101111111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11I_LC_14_5_2  (
            .in0(N__37979),
            .in1(N__35283),
            .in2(N__35239),
            .in3(N__35236),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_RNID11IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_5_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_22_c_inv_LC_14_5_5  (
            .in0(N__35080),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37977),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_14_5_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_14_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_23_c_inv_LC_14_5_7  (
            .in0(N__35211),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37978),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_14_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_14_6_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNIM1S01_12_LC_14_6_0  (
            .in0(N__37082),
            .in1(N__37950),
            .in2(N__35191),
            .in3(N__35152),
            .lcout(\current_shift_inst.PI_CTRL.error_control_RNIM1S01Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_14_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_14_6_1 .LUT_INIT=16'b0011111111001111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51J_LC_14_6_1  (
            .in0(N__35131),
            .in1(N__35079),
            .in2(N__37975),
            .in3(N__35062),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_RNII51JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_14_c_inv_LC_14_6_2  (
            .in0(N__35040),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37947),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_14_6_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_14_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_RNI1AJ_9_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35019),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_14_6_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_14_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_20_c_inv_LC_14_6_4  (
            .in0(N__38059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37949),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_14_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_14_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_inv_LC_14_6_6  (
            .in0(N__34983),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37948),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_14_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_14_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_26_c_inv_LC_14_7_1  (
            .in0(N__35514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37934),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_14_7_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_14_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_17_c_inv_LC_14_7_3  (
            .in0(N__35490),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37933),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_14_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_14_7_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_28_c_inv_LC_14_7_4  (
            .in0(N__37935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35470),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28 ),
            .ltout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_14_7_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_14_7_5 .LUT_INIT=16'b0011111111110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8J_LC_14_7_5  (
            .in0(N__35458),
            .in1(N__37936),
            .in2(N__35407),
            .in3(N__35404),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_27_c_RNILF8JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35382),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_14_8_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_14_8_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_21_c_inv_LC_14_8_2  (
            .in0(N__35339),
            .in1(N__37937),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_14_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_14_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI4JH5_16_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38004),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_14_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_14_8_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_24_c_inv_LC_14_8_4  (
            .in0(_gnd_net_),
            .in1(N__37938),
            .in2(_gnd_net_),
            .in3(N__35306),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_14_8_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_14_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI7MH5_19_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35651),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_14_8_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_14_8_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMI8D_9_LC_14_8_6  (
            .in0(N__38086),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_8_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_30_c_inv_LC_14_8_7  (
            .in0(N__37939),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35583),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_14_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_14_9_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0_9_LC_14_9_0  (
            .in0(N__41319),
            .in1(N__38467),
            .in2(_gnd_net_),
            .in3(N__35776),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a5_1_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_9_1 .LUT_INIT=16'b1101110111011100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_1_9_LC_14_9_1  (
            .in0(N__41594),
            .in1(N__41761),
            .in2(N__35563),
            .in3(N__38659),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_14_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_14_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_14_9_2 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_14_9_2  (
            .in0(N__41320),
            .in1(N__41596),
            .in2(N__35560),
            .in3(N__38429),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49939),
            .ce(N__36754),
            .sr(N__49421));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_14_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_14_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_14_9_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_14_9_5  (
            .in0(N__38468),
            .in1(N__41763),
            .in2(N__41630),
            .in3(N__38692),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49939),
            .ce(N__36754),
            .sr(N__49421));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_14_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_14_9_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_14_9_6  (
            .in0(N__41762),
            .in1(N__41595),
            .in2(_gnd_net_),
            .in3(N__41968),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49939),
            .ce(N__36754),
            .sr(N__49421));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_14_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_14_9_7 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_14_9_7  (
            .in0(N__35908),
            .in1(N__35922),
            .in2(N__36517),
            .in3(N__36477),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_14_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_14_10_1 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIR9HF91_12_LC_14_10_1  (
            .in0(N__41023),
            .in1(N__44053),
            .in2(N__40816),
            .in3(N__38524),
            .lcout(elapsed_time_ns_1_RNIR9HF91_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_10_2 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ8HF91_11_LC_14_10_2  (
            .in0(N__38548),
            .in1(N__44101),
            .in2(N__40818),
            .in3(N__41024),
            .lcout(elapsed_time_ns_1_RNIQ8HF91_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_10_3 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFJ2591_7_LC_14_10_3  (
            .in0(N__41025),
            .in1(N__35714),
            .in2(N__40817),
            .in3(N__47275),
            .lcout(elapsed_time_ns_1_RNIFJ2591_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_14_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_14_10_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_10_LC_14_10_4  (
            .in0(N__41444),
            .in1(N__38684),
            .in2(_gnd_net_),
            .in3(N__38469),
            .lcout(\phase_controller_inst1.stoper_tr.N_244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_14_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_14_10_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISAHF91_13_LC_14_10_7  (
            .in0(N__41022),
            .in1(N__44011),
            .in2(N__40815),
            .in3(N__38499),
            .lcout(elapsed_time_ns_1_RNISAHF91_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_11_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGK2591_8_LC_14_11_0  (
            .in0(N__35675),
            .in1(N__41054),
            .in2(N__47302),
            .in3(N__40822),
            .lcout(elapsed_time_ns_1_RNIGK2591_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_14_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_14_11_2 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_3_LC_14_11_2  (
            .in0(N__41770),
            .in1(N__38622),
            .in2(N__38643),
            .in3(N__41625),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_11_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIP7HF91_10_LC_14_11_3  (
            .in0(N__40821),
            .in1(N__38564),
            .in2(N__41061),
            .in3(N__43480),
            .lcout(elapsed_time_ns_1_RNIP7HF91_0_10),
            .ltout(elapsed_time_ns_1_RNIP7HF91_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_14_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_14_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_2_LC_14_11_4  (
            .in0(N__38494),
            .in1(N__38521),
            .in2(N__35722),
            .in3(N__38545),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_14_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_14_11_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_2_LC_14_11_5  (
            .in0(N__35707),
            .in1(N__40634),
            .in2(N__35686),
            .in3(N__35674),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_14_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_14_11_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_6_LC_14_11_6  (
            .in0(N__38470),
            .in1(_gnd_net_),
            .in2(N__35779),
            .in3(N__41624),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_14_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_14_11_7 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_0_2_LC_14_11_7  (
            .in0(N__38623),
            .in1(N__40685),
            .in2(N__38644),
            .in3(N__38608),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_12_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_9_LC_14_12_1  (
            .in0(N__38472),
            .in1(N__41310),
            .in2(_gnd_net_),
            .in3(N__41432),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_12_3 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_6_LC_14_12_3  (
            .in0(N__41433),
            .in1(N__41311),
            .in2(_gnd_net_),
            .in3(N__35772),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_12_4 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0_6_LC_14_12_4  (
            .in0(N__38683),
            .in1(N__38473),
            .in2(N__35761),
            .in3(N__41626),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_a2_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_12_5 .LUT_INIT=16'b1010101011111010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_0_1_LC_14_12_5  (
            .in0(N__41698),
            .in1(_gnd_net_),
            .in2(N__35758),
            .in3(N__38910),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_14_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_14_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_14_12_6 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_14_12_6  (
            .in0(N__38911),
            .in1(N__38896),
            .in2(N__35755),
            .in3(N__38849),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49921),
            .ce(N__36750),
            .sr(N__49439));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_14_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_14_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_14_12_7 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_14_12_7  (
            .in0(N__41699),
            .in1(N__38874),
            .in2(N__38856),
            .in3(N__38780),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49921),
            .ce(N__36750),
            .sr(N__49439));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_14_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_14_13_0 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL8GK01_19_LC_14_13_0  (
            .in0(N__45354),
            .in1(N__41875),
            .in2(N__41062),
            .in3(N__47173),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_14_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_14_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_14_13_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_14_13_2  (
            .in0(N__41751),
            .in1(N__41874),
            .in2(_gnd_net_),
            .in3(N__41629),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49916),
            .ce(N__36762),
            .sr(N__49450));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_13_3 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_13_3  (
            .in0(N__36420),
            .in1(N__35931),
            .in2(N__36448),
            .in3(N__35949),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_13_4 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_13_4  (
            .in0(N__35932),
            .in1(N__36447),
            .in2(N__35953),
            .in3(N__36421),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_13_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_14_13_5  (
            .in0(N__41627),
            .in1(N__41750),
            .in2(_gnd_net_),
            .in3(N__41503),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49916),
            .ce(N__36762),
            .sr(N__49450));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_14_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_14_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_14_13_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_14_13_6  (
            .in0(N__41749),
            .in1(N__41923),
            .in2(_gnd_net_),
            .in3(N__41628),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49916),
            .ce(N__36762),
            .sr(N__49450));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_14_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_14_13_7 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_14_13_7  (
            .in0(N__36478),
            .in1(N__35923),
            .in2(N__36516),
            .in3(N__35904),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_14_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_14_14_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_14_14_0  (
            .in0(N__35883),
            .in1(N__41197),
            .in2(N__46201),
            .in3(N__35843),
            .lcout(),
            .ltout(\phase_controller_inst2.start_timer_tr_RNO_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_14_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_14_14_1 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_14_14_1  (
            .in0(N__35817),
            .in1(N__36170),
            .in2(N__35797),
            .in3(N__44553),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49910),
            .ce(),
            .sr(N__49457));
    defparam \phase_controller_inst2.stoper_tr.running_LC_14_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_14_14_3 .LUT_INIT=16'b1000101011111010;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_14_14_3  (
            .in0(N__36190),
            .in1(N__35793),
            .in2(N__36142),
            .in3(N__36224),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49910),
            .ce(),
            .sr(N__49457));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_14_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_14_14_4 .LUT_INIT=16'b1101111111011101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIHOGI1_28_LC_14_14_4  (
            .in0(N__36223),
            .in1(N__37043),
            .in2(N__36795),
            .in3(N__36238),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_14_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36232),
            .in3(N__36125),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_14_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_14_6  (
            .in0(N__36222),
            .in1(N__36189),
            .in2(_gnd_net_),
            .in3(N__36163),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(\phase_controller_inst2.stoper_tr.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_14_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_14_14_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2_28_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36109),
            .in3(N__36099),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIQU8A2Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__36088),
            .in2(N__36082),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_15_1  (
            .in0(N__36743),
            .in1(N__36048),
            .in2(_gnd_net_),
            .in3(N__36034),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49906),
            .ce(),
            .sr(N__49464));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_15_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_15_2  (
            .in0(N__36747),
            .in1(N__36021),
            .in2(N__36031),
            .in3(N__36007),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49906),
            .ce(),
            .sr(N__49464));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_15_3  (
            .in0(N__36744),
            .in1(N__36003),
            .in2(_gnd_net_),
            .in3(N__35989),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49906),
            .ce(),
            .sr(N__49464));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_15_4  (
            .in0(N__36748),
            .in1(N__35985),
            .in2(_gnd_net_),
            .in3(N__35971),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49906),
            .ce(),
            .sr(N__49464));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_15_5  (
            .in0(N__36745),
            .in1(N__36387),
            .in2(_gnd_net_),
            .in3(N__36373),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49906),
            .ce(),
            .sr(N__49464));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_15_6  (
            .in0(N__36749),
            .in1(N__36369),
            .in2(_gnd_net_),
            .in3(N__36355),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49906),
            .ce(),
            .sr(N__49464));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_15_7  (
            .in0(N__36746),
            .in1(N__36351),
            .in2(_gnd_net_),
            .in3(N__36337),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49906),
            .ce(),
            .sr(N__49464));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_16_0  (
            .in0(N__36729),
            .in1(N__36333),
            .in2(_gnd_net_),
            .in3(N__36319),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49900),
            .ce(),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_16_1  (
            .in0(N__36696),
            .in1(N__36315),
            .in2(_gnd_net_),
            .in3(N__36301),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49900),
            .ce(),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_16_2  (
            .in0(N__36726),
            .in1(N__36291),
            .in2(_gnd_net_),
            .in3(N__36277),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49900),
            .ce(),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_16_3  (
            .in0(N__36697),
            .in1(N__36273),
            .in2(_gnd_net_),
            .in3(N__36259),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49900),
            .ce(),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_16_4  (
            .in0(N__36727),
            .in1(N__36255),
            .in2(_gnd_net_),
            .in3(N__36241),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49900),
            .ce(),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_16_5  (
            .in0(N__36698),
            .in1(N__36555),
            .in2(_gnd_net_),
            .in3(N__36541),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49900),
            .ce(),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_16_6  (
            .in0(N__36728),
            .in1(N__36534),
            .in2(_gnd_net_),
            .in3(N__36520),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49900),
            .ce(),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_16_7  (
            .in0(N__36699),
            .in1(N__36500),
            .in2(_gnd_net_),
            .in3(N__36481),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49900),
            .ce(),
            .sr(N__49471));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_17_0  (
            .in0(N__36692),
            .in1(N__36473),
            .in2(_gnd_net_),
            .in3(N__36451),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49895),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_17_1  (
            .in0(N__36722),
            .in1(N__36438),
            .in2(_gnd_net_),
            .in3(N__36424),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49895),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_17_2  (
            .in0(N__36693),
            .in1(N__36419),
            .in2(_gnd_net_),
            .in3(N__36403),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49895),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_17_3  (
            .in0(N__36723),
            .in1(N__36999),
            .in2(_gnd_net_),
            .in3(N__36400),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49895),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_17_4  (
            .in0(N__36694),
            .in1(N__37014),
            .in2(_gnd_net_),
            .in3(N__36397),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49895),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_17_5  (
            .in0(N__36724),
            .in1(N__36957),
            .in2(_gnd_net_),
            .in3(N__36394),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49895),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_17_6  (
            .in0(N__36695),
            .in1(N__36972),
            .in2(_gnd_net_),
            .in3(N__36853),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49895),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_17_7  (
            .in0(N__36725),
            .in1(N__36930),
            .in2(_gnd_net_),
            .in3(N__36850),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49895),
            .ce(),
            .sr(N__49480));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_18_0  (
            .in0(N__36688),
            .in1(N__36916),
            .in2(_gnd_net_),
            .in3(N__36847),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49889),
            .ce(),
            .sr(N__49487));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_18_1  (
            .in0(N__36719),
            .in1(N__36879),
            .in2(_gnd_net_),
            .in3(N__36844),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49889),
            .ce(),
            .sr(N__49487));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_18_2  (
            .in0(N__36689),
            .in1(N__36892),
            .in2(_gnd_net_),
            .in3(N__36841),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49889),
            .ce(),
            .sr(N__49487));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_18_3  (
            .in0(N__36720),
            .in1(N__36834),
            .in2(_gnd_net_),
            .in3(N__36820),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49889),
            .ce(),
            .sr(N__49487));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_18_4  (
            .in0(N__36690),
            .in1(N__36813),
            .in2(_gnd_net_),
            .in3(N__36799),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49889),
            .ce(),
            .sr(N__49487));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_18_5  (
            .in0(N__36721),
            .in1(N__36788),
            .in2(_gnd_net_),
            .in3(N__36766),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49889),
            .ce(),
            .sr(N__49487));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_18_6  (
            .in0(N__36691),
            .in1(N__37042),
            .in2(_gnd_net_),
            .in3(N__37060),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49889),
            .ce(),
            .sr(N__49487));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__48286),
            .in2(_gnd_net_),
            .in3(N__47968),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__47992),
            .in2(_gnd_net_),
            .in3(N__48013),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_14_19_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_14_19_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI1I3CP1_9_LC_14_19_2  (
            .in0(N__45208),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46023),
            .lcout(elapsed_time_ns_1_RNI1I3CP1_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_14_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_14_19_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4_2_LC_14_19_3  (
            .in0(N__42775),
            .in1(N__42646),
            .in2(_gnd_net_),
            .in3(N__39268),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_14_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_14_19_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_14_19_4  (
            .in0(N__37015),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37000),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__36973),
            .in2(_gnd_net_),
            .in3(N__36958),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_14_19_6  (
            .in0(N__36931),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36915),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_14_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_14_19_7 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_14_19_7  (
            .in0(N__36891),
            .in1(_gnd_net_),
            .in2(N__36880),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_14_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_14_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_14_20_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_14_20_1  (
            .in0(N__47106),
            .in1(N__38322),
            .in2(_gnd_net_),
            .in3(N__42205),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49875),
            .ce(N__49121),
            .sr(N__49502));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_14_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_14_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_14_20_5 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_14_20_5  (
            .in0(N__47107),
            .in1(N__45757),
            .in2(N__45602),
            .in3(N__46826),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49875),
            .ce(N__49121),
            .sr(N__49502));
    defparam \phase_controller_inst1.state_2_LC_14_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_14_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_14_22_6 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst1.state_2_LC_14_22_6  (
            .in0(N__38294),
            .in1(N__46587),
            .in2(N__44640),
            .in3(N__38255),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49865),
            .ce(),
            .sr(N__49514));
    defparam \phase_controller_inst1.T01_LC_14_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_14_23_0 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst1.T01_LC_14_23_0  (
            .in0(N__38202),
            .in1(N__38256),
            .in2(_gnd_net_),
            .in3(N__46588),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49860),
            .ce(),
            .sr(N__49518));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_15_5_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_15_5_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_15_5_0 .LUT_INIT=16'b0100010011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_15_5_0  (
            .in0(N__37713),
            .in1(N__37498),
            .in2(N__37326),
            .in3(N__38191),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49965),
            .ce(),
            .sr(N__49406));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2 .LUT_INIT=16'b0000000111110101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_15_6_2  (
            .in0(N__37501),
            .in1(N__37284),
            .in2(N__37714),
            .in3(N__38122),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49960),
            .ce(),
            .sr(N__49408));
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_15_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_15_6_6 .LUT_INIT=16'b0101111110101111;
    LogicCell40 \current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6I_LC_15_6_6  (
            .in0(N__38058),
            .in1(N__38035),
            .in2(N__37984),
            .in3(N__37738),
            .lcout(\current_shift_inst.PI_CTRL.un7_integrator_1_cry_19_c_RNING6IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_15_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_15_7_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_15_7_4 .LUT_INIT=16'b0000000110111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_15_7_4  (
            .in0(N__37709),
            .in1(N__37497),
            .in2(N__37327),
            .in3(N__37123),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49954),
            .ce(),
            .sr(N__49410));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_8_0 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVEIF91_25_LC_15_8_0  (
            .in0(N__40972),
            .in1(N__38374),
            .in2(N__44206),
            .in3(N__40779),
            .lcout(elapsed_time_ns_1_RNIVEIF91_0_25),
            .ltout(elapsed_time_ns_1_RNIVEIF91_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_6_15_LC_15_8_1  (
            .in0(N__38364),
            .in1(N__38352),
            .in2(N__38368),
            .in3(N__38583),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_6Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_8_4 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2IIF91_28_LC_15_8_4  (
            .in0(N__40973),
            .in1(N__38365),
            .in2(N__44857),
            .in3(N__40780),
            .lcout(elapsed_time_ns_1_RNI2IIF91_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_15_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_15_8_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1HIF91_27_LC_15_8_6  (
            .in0(N__40974),
            .in1(N__44914),
            .in2(N__38356),
            .in3(N__40781),
            .lcout(elapsed_time_ns_1_RNI1HIF91_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_15_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_15_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_15_LC_15_9_0  (
            .in0(N__40255),
            .in1(N__38344),
            .in2(N__40597),
            .in3(N__38331),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_19_LC_15_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_19_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_19_LC_15_9_2 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIB51JG_19_LC_15_9_2  (
            .in0(N__49580),
            .in1(N__41173),
            .in2(N__47455),
            .in3(N__45290),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_9_3 .LUT_INIT=16'b1111100011111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJ_31_LC_15_9_3  (
            .in0(N__44695),
            .in1(N__49581),
            .in2(N__38338),
            .in3(N__47719),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK4GOJZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_9_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRAIF91_21_LC_15_9_4  (
            .in0(N__44377),
            .in1(N__41007),
            .in2(N__38335),
            .in3(N__40279),
            .lcout(elapsed_time_ns_1_RNIRAIF91_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_9_5 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISBIF91_22_LC_15_9_5  (
            .in0(N__38332),
            .in1(N__44338),
            .in2(N__41049),
            .in3(N__40785),
            .lcout(elapsed_time_ns_1_RNISBIF91_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_9_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFON8L_31_LC_15_9_6  (
            .in0(N__41395),
            .in1(N__44694),
            .in2(_gnd_net_),
            .in3(N__41380),
            .lcout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i ),
            .ltout(\delay_measurement_inst.delay_tr_timer.un4_elapsed_time_tr_1_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_15_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_15_9_7 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0GIF91_26_LC_15_9_7  (
            .in0(N__38584),
            .in1(N__44161),
            .in2(N__38587),
            .in3(N__40784),
            .lcout(elapsed_time_ns_1_RNI0GIF91_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_15_10_0 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_15_10_0  (
            .in0(N__41775),
            .in1(N__41448),
            .in2(N__41623),
            .in3(N__38419),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(N__50322),
            .sr(N__49422));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_15_10_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_15_10_1  (
            .in0(N__38414),
            .in1(N__41568),
            .in2(N__38571),
            .in3(N__41771),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(N__50322),
            .sr(N__49422));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_15_10_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_15_10_2  (
            .in0(N__41772),
            .in1(N__38417),
            .in2(N__41621),
            .in3(N__38546),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(N__50322),
            .sr(N__49422));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_15_10_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_15_10_3  (
            .in0(N__38415),
            .in1(N__38523),
            .in2(N__41632),
            .in3(N__41773),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(N__50322),
            .sr(N__49422));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_15_10_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_15_10_4  (
            .in0(N__41774),
            .in1(N__38418),
            .in2(N__41622),
            .in3(N__38495),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(N__50322),
            .sr(N__49422));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_10_5 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUCHF91_15_LC_15_10_5  (
            .in0(N__43930),
            .in1(N__38471),
            .in2(N__41050),
            .in3(N__40788),
            .lcout(elapsed_time_ns_1_RNIUCHF91_0_15),
            .ltout(elapsed_time_ns_1_RNIUCHF91_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_15_10_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_15_10_6  (
            .in0(N__41776),
            .in1(N__41600),
            .in2(N__38434),
            .in3(N__38688),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(N__50322),
            .sr(N__49422));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_15_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_15_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_15_10_7 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_15_10_7  (
            .in0(N__38416),
            .in1(N__41317),
            .in2(N__41631),
            .in3(N__38380),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49940),
            .ce(N__50322),
            .sr(N__49422));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_15_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_15_11_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_9_LC_15_11_0  (
            .in0(N__41955),
            .in1(N__41911),
            .in2(N__41498),
            .in3(N__41861),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_i_o2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_15_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_15_11_1 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAE2591_2_LC_15_11_1  (
            .in0(N__38607),
            .in1(N__41055),
            .in2(N__47368),
            .in3(N__40819),
            .lcout(elapsed_time_ns_1_RNIAE2591_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_7_LC_15_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_7_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_7_LC_15_11_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITAPC7_7_LC_15_11_2  (
            .in0(N__40856),
            .in1(N__41168),
            .in2(_gnd_net_),
            .in3(N__40835),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_386_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_15_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_15_11_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIEC3FA_1_LC_15_11_3  (
            .in0(N__47311),
            .in1(_gnd_net_),
            .in2(N__38662),
            .in3(N__47711),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_15_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_15_11_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_2_LC_15_11_4  (
            .in0(N__41956),
            .in1(N__41068),
            .in2(N__41918),
            .in3(N__38655),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2 ),
            .ltout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_15_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_15_11_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5_1_LC_15_11_5  (
            .in0(N__38593),
            .in1(N__41593),
            .in2(N__38626),
            .in3(N__38621),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_a5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_11_6 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2_1_LC_15_11_6  (
            .in0(N__40674),
            .in1(N__38606),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_f0_0_o2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_19_LC_15_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_19_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_19_LC_15_11_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8S8BA_19_LC_15_11_7  (
            .in0(N__41169),
            .in1(N__40857),
            .in2(N__40840),
            .in3(N__47451),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_12_0 .LUT_INIT=16'b1011111110101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIS41A01_1_LC_15_12_0  (
            .in0(N__45348),
            .in1(N__41056),
            .in2(N__47332),
            .in3(N__38909),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_15_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_15_12_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII6NQL1_1_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38914),
            .in3(N__41365),
            .lcout(elapsed_time_ns_1_RNII6NQL1_0_1),
            .ltout(elapsed_time_ns_1_RNII6NQL1_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_15_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_15_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_15_12_2 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_15_12_2  (
            .in0(N__38895),
            .in1(N__38839),
            .in2(N__38884),
            .in3(N__38881),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49927),
            .ce(N__50323),
            .sr(N__49433));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_15_12_3 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_15_12_3  (
            .in0(N__38838),
            .in1(N__41769),
            .in2(N__38790),
            .in3(N__40630),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49927),
            .ce(N__50323),
            .sr(N__49433));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_12_4 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISCJF91_31_LC_15_12_4  (
            .in0(N__41764),
            .in1(N__44693),
            .in2(N__41060),
            .in3(N__40820),
            .lcout(elapsed_time_ns_1_RNISCJF91_0_31),
            .ltout(elapsed_time_ns_1_RNISCJF91_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_15_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_15_12_5 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_15_12_5  (
            .in0(N__38837),
            .in1(N__38875),
            .in2(N__38863),
            .in3(N__38781),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49927),
            .ce(N__50323),
            .sr(N__49433));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_15_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_15_12_6 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_15_12_6  (
            .in0(N__41100),
            .in1(N__38772),
            .in2(N__41802),
            .in3(N__38843),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49927),
            .ce(N__50323),
            .sr(N__49433));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_15_12_7 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_15_12_7  (
            .in0(N__41138),
            .in1(N__41768),
            .in2(N__38855),
            .in3(N__38782),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49927),
            .ce(N__50323),
            .sr(N__49433));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__38713),
            .in2(N__38722),
            .in3(N__47669),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__38698),
            .in2(N__38707),
            .in3(N__47656),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_15_13_2  (
            .in0(N__47623),
            .in1(N__39061),
            .in2(N__39049),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_13_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_15_13_3  (
            .in0(N__47605),
            .in1(N__39040),
            .in2(N__39034),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__39025),
            .in2(N__39019),
            .in3(N__47584),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__39010),
            .in2(N__39004),
            .in3(N__47566),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__38992),
            .in2(N__38980),
            .in3(N__47548),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_15_13_7  (
            .in0(N__47527),
            .in1(N__38971),
            .in2(N__38959),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__38950),
            .in2(N__38941),
            .in3(N__47941),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__38932),
            .in2(N__38923),
            .in3(N__47923),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_14_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_15_14_2  (
            .in0(N__47905),
            .in1(N__39142),
            .in2(N__39154),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__39136),
            .in2(N__39127),
            .in3(N__47887),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__39118),
            .in2(N__39109),
            .in3(N__47869),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__39100),
            .in2(N__39091),
            .in3(N__47851),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__39079),
            .in2(N__39070),
            .in3(N__47833),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__41974),
            .in2(N__41989),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_15_15_0  (
            .in0(_gnd_net_),
            .in1(N__41815),
            .in2(N__41839),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_15_15_1  (
            .in0(_gnd_net_),
            .in1(N__48847),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(N__39196),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__39184),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__45025),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(N__45037),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__44953),
            .in2(N__48178),
            .in3(N__39172),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39169),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_15_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_15_16_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_7_15_LC_15_16_0  (
            .in0(N__42045),
            .in1(N__39249),
            .in2(N__39166),
            .in3(N__39258),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_7Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_15_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_15_16_1 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4HV8E1_30_LC_15_16_1  (
            .in0(N__45861),
            .in1(N__39489),
            .in2(N__45511),
            .in3(N__39165),
            .lcout(elapsed_time_ns_1_RNI4HV8E1_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_15_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_15_16_2 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI8KU8E1_25_LC_15_16_2  (
            .in0(N__45459),
            .in1(N__45868),
            .in2(N__42475),
            .in3(N__45169),
            .lcout(elapsed_time_ns_1_RNI8KU8E1_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_15_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_15_16_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNILGKEE1_4_LC_15_16_3  (
            .in0(N__45860),
            .in1(N__45455),
            .in2(N__39296),
            .in3(N__39219),
            .lcout(elapsed_time_ns_1_RNILGKEE1_0_4),
            .ltout(elapsed_time_ns_1_RNILGKEE1_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_15_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_15_16_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3_2_LC_15_16_4  (
            .in0(N__42302),
            .in1(N__42954),
            .in2(N__39271),
            .in3(N__43375),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_1_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_15_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_15_16_5 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4GU8E1_21_LC_15_16_5  (
            .in0(N__39259),
            .in1(N__42034),
            .in2(N__45905),
            .in3(N__45458),
            .lcout(elapsed_time_ns_1_RNI4GU8E1_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_15_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_15_16_6 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2DT8E1_10_LC_15_16_6  (
            .in0(N__45456),
            .in1(N__43297),
            .in2(N__45927),
            .in3(N__39339),
            .lcout(elapsed_time_ns_1_RNI2DT8E1_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_15_16_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_15_16_7 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNICOU8E1_29_LC_15_16_7  (
            .in0(N__39250),
            .in1(N__39517),
            .in2(N__45904),
            .in3(N__45457),
            .lcout(elapsed_time_ns_1_RNICOU8E1_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_17_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__39723),
            .in2(N__39430),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49901),
            .ce(N__39451),
            .sr(N__49472));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__39702),
            .in2(N__39760),
            .in3(N__39205),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49901),
            .ce(N__39451),
            .sr(N__49472));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__39724),
            .in2(N__39679),
            .in3(N__39202),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49901),
            .ce(N__39451),
            .sr(N__49472));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__39703),
            .in2(N__39651),
            .in3(N__39199),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49901),
            .ce(N__39451),
            .sr(N__49472));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__39678),
            .in2(N__39621),
            .in3(N__39361),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49901),
            .ce(N__39451),
            .sr(N__49472));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__39588),
            .in2(N__39652),
            .in3(N__39346),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49901),
            .ce(N__39451),
            .sr(N__49472));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__39555),
            .in2(N__39622),
            .in3(N__39343),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49901),
            .ce(N__39451),
            .sr(N__49472));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__39987),
            .in2(N__39592),
            .in3(N__39325),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49901),
            .ce(N__39451),
            .sr(N__49472));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__39960),
            .in2(N__39562),
            .in3(N__39322),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49896),
            .ce(N__39450),
            .sr(N__49481));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__39936),
            .in2(N__39991),
            .in3(N__39319),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49896),
            .ce(N__39450),
            .sr(N__49481));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__39961),
            .in2(N__39912),
            .in3(N__39316),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49896),
            .ce(N__39450),
            .sr(N__49481));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__39937),
            .in2(N__39882),
            .in3(N__39313),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49896),
            .ce(N__39450),
            .sr(N__49481));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__39849),
            .in2(N__39913),
            .in3(N__39310),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49896),
            .ce(N__39450),
            .sr(N__49481));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_18_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__39819),
            .in2(N__39883),
            .in3(N__39400),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49896),
            .ce(N__39450),
            .sr(N__49481));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_18_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_18_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__39789),
            .in2(N__39853),
            .in3(N__39397),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49896),
            .ce(N__39450),
            .sr(N__49481));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_18_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_18_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__40239),
            .in2(N__39823),
            .in3(N__39394),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49896),
            .ce(N__39450),
            .sr(N__49481));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_19_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_19_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__40209),
            .in2(N__39793),
            .in3(N__39391),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49890),
            .ce(N__39449),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_19_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_19_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__40243),
            .in2(N__40182),
            .in3(N__39388),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49890),
            .ce(N__39449),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_19_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_19_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__40155),
            .in2(N__40213),
            .in3(N__39385),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49890),
            .ce(N__39449),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_19_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_19_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__40131),
            .in2(N__40183),
            .in3(N__39382),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49890),
            .ce(N__39449),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_19_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_19_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__40156),
            .in2(N__40107),
            .in3(N__39379),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49890),
            .ce(N__39449),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_19_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_19_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__40077),
            .in2(N__40135),
            .in3(N__39376),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49890),
            .ce(N__39449),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_19_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_19_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__40050),
            .in2(N__40108),
            .in3(N__39529),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49890),
            .ce(N__39449),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_19_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_19_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__40078),
            .in2(N__40023),
            .in3(N__39526),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49890),
            .ce(N__39449),
            .sr(N__49488));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_20_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_20_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__40551),
            .in2(N__40057),
            .in3(N__39523),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49882),
            .ce(N__39448),
            .sr(N__49493));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_20_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_20_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__40024),
            .in2(N__40530),
            .in3(N__39520),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49882),
            .ce(N__39448),
            .sr(N__49493));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_20_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__40552),
            .in2(N__40504),
            .in3(N__39496),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49882),
            .ce(N__39448),
            .sr(N__49493));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_20_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__40342),
            .in2(N__40531),
            .in3(N__39469),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49882),
            .ce(N__39448),
            .sr(N__49493));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_20_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_20_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39466),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49882),
            .ce(N__39448),
            .sr(N__49493));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_20_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_20_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39423),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49882),
            .ce(N__39448),
            .sr(N__49493));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_21_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_21_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_15_21_0  (
            .in0(N__40476),
            .in1(N__39422),
            .in2(_gnd_net_),
            .in3(N__39403),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__49876),
            .ce(N__40318),
            .sr(N__49503));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_21_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_21_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_15_21_1  (
            .in0(N__40480),
            .in1(N__39746),
            .in2(_gnd_net_),
            .in3(N__39727),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__49876),
            .ce(N__40318),
            .sr(N__49503));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_21_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_15_21_2  (
            .in0(N__40477),
            .in1(N__39722),
            .in2(_gnd_net_),
            .in3(N__39706),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__49876),
            .ce(N__40318),
            .sr(N__49503));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_21_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_15_21_3  (
            .in0(N__40481),
            .in1(N__39696),
            .in2(_gnd_net_),
            .in3(N__39682),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__49876),
            .ce(N__40318),
            .sr(N__49503));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_21_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_21_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_15_21_4  (
            .in0(N__40478),
            .in1(N__39674),
            .in2(_gnd_net_),
            .in3(N__39655),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__49876),
            .ce(N__40318),
            .sr(N__49503));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_21_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_21_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_15_21_5  (
            .in0(N__40482),
            .in1(N__39639),
            .in2(_gnd_net_),
            .in3(N__39625),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__49876),
            .ce(N__40318),
            .sr(N__49503));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_21_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_21_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_15_21_6  (
            .in0(N__40479),
            .in1(N__39609),
            .in2(_gnd_net_),
            .in3(N__39595),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__49876),
            .ce(N__40318),
            .sr(N__49503));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_21_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_21_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_15_21_7  (
            .in0(N__40483),
            .in1(N__39581),
            .in2(_gnd_net_),
            .in3(N__39565),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__49876),
            .ce(N__40318),
            .sr(N__49503));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_22_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_15_22_0  (
            .in0(N__40404),
            .in1(N__39554),
            .in2(_gnd_net_),
            .in3(N__39532),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_22_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__49870),
            .ce(N__40326),
            .sr(N__49508));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_22_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_22_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_15_22_1  (
            .in0(N__40443),
            .in1(N__39980),
            .in2(_gnd_net_),
            .in3(N__39964),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__49870),
            .ce(N__40326),
            .sr(N__49508));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_22_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_15_22_2  (
            .in0(N__40401),
            .in1(N__39954),
            .in2(_gnd_net_),
            .in3(N__39940),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__49870),
            .ce(N__40326),
            .sr(N__49508));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_22_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_15_22_3  (
            .in0(N__40440),
            .in1(N__39930),
            .in2(_gnd_net_),
            .in3(N__39916),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__49870),
            .ce(N__40326),
            .sr(N__49508));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_22_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_15_22_4  (
            .in0(N__40402),
            .in1(N__39900),
            .in2(_gnd_net_),
            .in3(N__39886),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__49870),
            .ce(N__40326),
            .sr(N__49508));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_22_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_22_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_15_22_5  (
            .in0(N__40441),
            .in1(N__39870),
            .in2(_gnd_net_),
            .in3(N__39856),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__49870),
            .ce(N__40326),
            .sr(N__49508));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_22_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_22_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_15_22_6  (
            .in0(N__40403),
            .in1(N__39842),
            .in2(_gnd_net_),
            .in3(N__39826),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__49870),
            .ce(N__40326),
            .sr(N__49508));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_22_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_22_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_15_22_7  (
            .in0(N__40442),
            .in1(N__39812),
            .in2(_gnd_net_),
            .in3(N__39796),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__49870),
            .ce(N__40326),
            .sr(N__49508));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_23_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_23_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_23_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_15_23_0  (
            .in0(N__40457),
            .in1(N__39782),
            .in2(_gnd_net_),
            .in3(N__39763),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_15_23_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__49866),
            .ce(N__40325),
            .sr(N__49515));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_23_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_23_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_23_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_15_23_1  (
            .in0(N__40453),
            .in1(N__40238),
            .in2(_gnd_net_),
            .in3(N__40216),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__49866),
            .ce(N__40325),
            .sr(N__49515));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_23_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_23_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_23_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_15_23_2  (
            .in0(N__40458),
            .in1(N__40202),
            .in2(_gnd_net_),
            .in3(N__40186),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__49866),
            .ce(N__40325),
            .sr(N__49515));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_23_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_23_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_15_23_3  (
            .in0(N__40454),
            .in1(N__40175),
            .in2(_gnd_net_),
            .in3(N__40159),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__49866),
            .ce(N__40325),
            .sr(N__49515));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_23_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_23_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_23_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_15_23_4  (
            .in0(N__40459),
            .in1(N__40154),
            .in2(_gnd_net_),
            .in3(N__40138),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__49866),
            .ce(N__40325),
            .sr(N__49515));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_23_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_23_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_15_23_5  (
            .in0(N__40455),
            .in1(N__40130),
            .in2(_gnd_net_),
            .in3(N__40111),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__49866),
            .ce(N__40325),
            .sr(N__49515));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_23_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_23_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_15_23_6  (
            .in0(N__40460),
            .in1(N__40095),
            .in2(_gnd_net_),
            .in3(N__40081),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__49866),
            .ce(N__40325),
            .sr(N__49515));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_23_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_23_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_23_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_15_23_7  (
            .in0(N__40456),
            .in1(N__40076),
            .in2(_gnd_net_),
            .in3(N__40060),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__49866),
            .ce(N__40325),
            .sr(N__49515));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_24_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_15_24_0  (
            .in0(N__40461),
            .in1(N__40049),
            .in2(_gnd_net_),
            .in3(N__40027),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_15_24_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__49861),
            .ce(N__40327),
            .sr(N__49519));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_24_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_24_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_15_24_1  (
            .in0(N__40465),
            .in1(N__40016),
            .in2(_gnd_net_),
            .in3(N__39994),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__49861),
            .ce(N__40327),
            .sr(N__49519));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_24_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_24_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_15_24_2  (
            .in0(N__40462),
            .in1(N__40550),
            .in2(_gnd_net_),
            .in3(N__40534),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__49861),
            .ce(N__40327),
            .sr(N__49519));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_24_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_15_24_3  (
            .in0(N__40466),
            .in1(N__40523),
            .in2(_gnd_net_),
            .in3(N__40507),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__49861),
            .ce(N__40327),
            .sr(N__49519));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_24_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_15_24_4  (
            .in0(N__40463),
            .in1(N__40500),
            .in2(_gnd_net_),
            .in3(N__40486),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__49861),
            .ce(N__40327),
            .sr(N__49519));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_24_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_24_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_24_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_15_24_5  (
            .in0(N__40341),
            .in1(N__40464),
            .in2(_gnd_net_),
            .in3(N__40345),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49861),
            .ce(N__40327),
            .sr(N__49519));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_16_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_16_8_2 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3JIF91_29_LC_16_8_2  (
            .in0(N__40264),
            .in1(N__44785),
            .in2(N__41031),
            .in3(N__40778),
            .lcout(elapsed_time_ns_1_RNI3JIF91_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_16_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_16_8_4 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQ9IF91_20_LC_16_8_4  (
            .in0(N__44416),
            .in1(N__40285),
            .in2(N__41029),
            .in3(N__40776),
            .lcout(elapsed_time_ns_1_RNIQ9IF91_0_20),
            .ltout(elapsed_time_ns_1_RNIQ9IF91_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_8_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_7_15_LC_16_8_5  (
            .in0(N__40278),
            .in1(N__40563),
            .in2(N__40267),
            .in3(N__40263),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_7Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_8_6 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNITCIF91_23_LC_16_8_6  (
            .in0(N__44293),
            .in1(N__40249),
            .in2(N__41030),
            .in3(N__40777),
            .lcout(elapsed_time_ns_1_RNITCIF91_0_23),
            .ltout(elapsed_time_ns_1_RNITCIF91_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_16_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_16_8_7 .LUT_INIT=16'b1111110011111100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_15_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__40584),
            .in2(N__40600),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_o5_0_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_9_0 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUDIF91_24_LC_16_9_0  (
            .in0(N__41033),
            .in1(N__44248),
            .in2(N__40588),
            .in3(N__40783),
            .lcout(elapsed_time_ns_1_RNIUDIF91_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_16_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_16_9_1 .LUT_INIT=16'b0011001000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3GEH5_15_LC_16_9_1  (
            .in0(N__43929),
            .in1(N__47152),
            .in2(N__47776),
            .in3(N__40705),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_9_2 .LUT_INIT=16'b0101010101010001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_16_9_2  (
            .in0(N__44680),
            .in1(N__40861),
            .in2(N__40573),
            .in3(N__40839),
            .lcout(\delay_measurement_inst.delay_tr9 ),
            .ltout(\delay_measurement_inst.delay_tr9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_16_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_16_9_3 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1A1A01_6_LC_16_9_3  (
            .in0(N__47743),
            .in1(N__40638),
            .in2(N__40570),
            .in3(N__41034),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_9_6 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG3GK01_14_LC_16_9_6  (
            .in0(N__41035),
            .in1(N__41443),
            .in2(N__45334),
            .in3(N__47775),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_16_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_16_9_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRBJF91_30_LC_16_9_7  (
            .in0(N__40782),
            .in1(N__41032),
            .in2(N__40567),
            .in3(N__44722),
            .lcout(elapsed_time_ns_1_RNIRBJF91_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_16_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_16_10_0 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK7GK01_18_LC_16_10_0  (
            .in0(N__41039),
            .in1(N__41488),
            .in2(N__45332),
            .in3(N__47233),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_16_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_16_10_1 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4D1A01_9_LC_16_10_1  (
            .in0(N__41318),
            .in1(N__47794),
            .in2(N__45335),
            .in3(N__41042),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_10_2 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICG2591_4_LC_16_10_2  (
            .in0(N__41040),
            .in1(N__41096),
            .in2(N__47410),
            .in3(N__40787),
            .lcout(elapsed_time_ns_1_RNICG2591_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJL0B1_24_LC_16_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJL0B1_24_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJL0B1_24_LC_16_10_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJL0B1_24_LC_16_10_3  (
            .in0(N__44721),
            .in1(N__44784),
            .in2(_gnd_net_),
            .in3(N__44244),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_23_LC_16_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_23_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_23_LC_16_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQVV04_23_LC_16_10_4  (
            .in0(N__44289),
            .in1(N__44157),
            .in2(N__40843),
            .in3(N__40870),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_16_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_16_10_5 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDH2591_5_LC_16_10_5  (
            .in0(N__40786),
            .in1(N__47422),
            .in2(N__41139),
            .in3(N__41041),
            .lcout(elapsed_time_ns_1_RNIDH2591_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_10_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIO7LR2_9_LC_16_10_6  (
            .in0(N__47793),
            .in1(N__40606),
            .in2(_gnd_net_),
            .in3(N__47245),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_16_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_16_10_7 .LUT_INIT=16'b1111101011111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII5GK01_16_LC_16_10_7  (
            .in0(N__47212),
            .in1(N__41963),
            .in2(N__45336),
            .in3(N__41043),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_16_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_16_11_0 .LUT_INIT=16'b1111110011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC8TA1_3_LC_16_11_0  (
            .in0(N__40684),
            .in1(N__41361),
            .in2(N__47386),
            .in3(N__41045),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_16_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_16_11_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIK8NQL1_3_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40699),
            .in3(N__45333),
            .lcout(elapsed_time_ns_1_RNIK8NQL1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_16_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_16_11_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINBNQL1_6_LC_16_11_2  (
            .in0(N__40651),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41359),
            .lcout(elapsed_time_ns_1_RNINBNQL1_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIUG5P1_10_LC_16_11_3  (
            .in0(N__44094),
            .in1(N__44046),
            .in2(N__44007),
            .in3(N__43476),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_353 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_353_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIE4F2_7_LC_16_11_4  (
            .in0(N__43916),
            .in1(N__47292),
            .in2(N__41176),
            .in3(N__47265),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_382 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_11_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8765M1_16_LC_16_11_5  (
            .in0(N__41360),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41155),
            .lcout(elapsed_time_ns_1_RNI8765M1_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_11_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIA965M1_18_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(N__41358),
            .in2(_gnd_net_),
            .in3(N__41149),
            .lcout(elapsed_time_ns_1_RNIA965M1_0_18),
            .ltout(elapsed_time_ns_1_RNIA965M1_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_11_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3_2_LC_16_11_7  (
            .in0(N__41860),
            .in1(N__41125),
            .in2(N__41107),
            .in3(N__41089),
            .lcout(\phase_controller_inst1.stoper_tr.target_time_4_i_a2_1_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_12_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI9865M1_17_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__40888),
            .in2(_gnd_net_),
            .in3(N__41362),
            .lcout(elapsed_time_ns_1_RNI9865M1_0_17),
            .ltout(elapsed_time_ns_1_RNI9865M1_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_12_1 .LUT_INIT=16'b1111111110111000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ6GK01_17_LC_16_12_1  (
            .in0(N__47193),
            .in1(N__41044),
            .in2(N__40891),
            .in3(N__45314),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_latch_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_16_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_16_12_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBA65M1_19_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__40882),
            .in2(_gnd_net_),
            .in3(N__41364),
            .lcout(elapsed_time_ns_1_RNIBA65M1_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG7AP1_20_LC_16_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG7AP1_20_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG7AP1_20_LC_16_12_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIG7AP1_20_LC_16_12_3  (
            .in0(N__44907),
            .in1(N__44196),
            .in2(N__44853),
            .in3(N__44409),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto31_0_o2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_16_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_16_12_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHSKS_21_LC_16_12_4  (
            .in0(N__44331),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44370),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lt31_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_12_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6565M1_14_LC_16_12_5  (
            .in0(N__41363),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41458),
            .lcout(elapsed_time_ns_1_RNI6565M1_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_12_6 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM1MGL_31_LC_16_12_6  (
            .in0(N__49582),
            .in1(N__41391),
            .in2(N__44692),
            .in3(N__41376),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_16_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_16_12_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIQENQL1_9_LC_16_12_7  (
            .in0(N__41332),
            .in1(_gnd_net_),
            .in2(N__41323),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNIQENQL1_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_13_0 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_16_13_0  (
            .in0(N__50292),
            .in1(N__45184),
            .in2(N__50038),
            .in3(N__47679),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__41262),
            .in2(_gnd_net_),
            .in3(N__41222),
            .lcout(),
            .ltout(\phase_controller_inst2.start_timer_hc_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_hc_LC_16_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_16_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_16_13_2 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_16_13_2  (
            .in0(N__44552),
            .in1(N__41274),
            .in2(N__41281),
            .in3(N__46152),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_13_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__46135),
            .in2(_gnd_net_),
            .in3(N__46151),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_16_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_16_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNIG7JF_2_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__41189),
            .in2(_gnd_net_),
            .in3(N__46190),
            .lcout(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_2_LC_16_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_16_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_16_13_7 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst2.state_2_LC_16_13_7  (
            .in0(N__41190),
            .in1(N__41263),
            .in2(N__46197),
            .in3(N__41223),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49928),
            .ce(),
            .sr(N__49434));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_14_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_16_14_0  (
            .in0(N__47814),
            .in1(N__48093),
            .in2(N__41887),
            .in3(N__41932),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_14_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_16_14_1  (
            .in0(N__41931),
            .in1(N__47815),
            .in2(N__48097),
            .in3(N__41883),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_16_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_16_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_16_14_2 .LUT_INIT=16'b0011001000110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_16_14_2  (
            .in0(N__41967),
            .in1(N__41798),
            .in2(N__41655),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49922),
            .ce(N__50320),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_16_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_16_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_16_14_3 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_16_14_3  (
            .in0(N__41799),
            .in1(N__41922),
            .in2(_gnd_net_),
            .in3(N__41647),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49922),
            .ce(N__50320),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_16_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_16_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_16_14_4 .LUT_INIT=16'b0011001000110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_16_14_4  (
            .in0(N__41868),
            .in1(N__41801),
            .in2(N__41656),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49922),
            .ce(N__50320),
            .sr(N__49440));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_14_5 .LUT_INIT=16'b1101111100001101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_16_14_5  (
            .in0(N__48069),
            .in1(N__41467),
            .in2(N__48046),
            .in3(N__41823),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_14_6 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_16_14_6  (
            .in0(N__41466),
            .in1(N__48042),
            .in2(N__41827),
            .in3(N__48070),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_16_14_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_16_14_7  (
            .in0(N__41800),
            .in1(N__41648),
            .in2(_gnd_net_),
            .in3(N__41502),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49922),
            .ce(N__50320),
            .sr(N__49440));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_16_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_16_15_0 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3ET8E1_11_LC_16_15_0  (
            .in0(N__42382),
            .in1(N__45903),
            .in2(N__43259),
            .in3(N__45466),
            .lcout(elapsed_time_ns_1_RNI3ET8E1_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_16_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_16_15_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_31_LC_16_15_1  (
            .in0(N__45311),
            .in1(N__49584),
            .in2(_gnd_net_),
            .in3(N__42363),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4NZ0Z_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_16_15_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_16_15_2 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4FT8E1_12_LC_16_15_2  (
            .in0(N__42400),
            .in1(N__43208),
            .in2(N__42100),
            .in3(N__45465),
            .lcout(elapsed_time_ns_1_RNI4FT8E1_0_12),
            .ltout(elapsed_time_ns_1_RNI4FT8E1_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_16_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_16_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_2_2_LC_16_15_3  (
            .in0(N__44971),
            .in1(N__43249),
            .in2(N__42097),
            .in3(N__43298),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_a2_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_16_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_16_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPR8P8_10_LC_16_15_4  (
            .in0(N__42094),
            .in1(N__42082),
            .in2(N__42070),
            .in3(N__45043),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlt31_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_16_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_16_15_5 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIP0VUB_31_LC_16_15_5  (
            .in0(N__44664),
            .in1(N__42135),
            .in2(N__42055),
            .in3(N__47718),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_369 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_16_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_16_15_6 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI0TDSM_31_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42052),
            .in3(N__45312),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_367_clk ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_367_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_16_15_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_16_15_7 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI3FU8E1_20_LC_16_15_7  (
            .in0(N__45902),
            .in1(N__42015),
            .in2(N__42049),
            .in3(N__42046),
            .lcout(elapsed_time_ns_1_RNI3FU8E1_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_16_16_0  (
            .in0(N__42345),
            .in1(N__42033),
            .in2(N__42016),
            .in3(N__42117),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_16_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_16_16_1 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5HU8E1_22_LC_16_16_1  (
            .in0(N__45463),
            .in1(N__42346),
            .in2(N__42454),
            .in3(N__45874),
            .lcout(elapsed_time_ns_1_RNI5HU8E1_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_16_16_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_16_16_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI6IU8E1_23_LC_16_16_2  (
            .in0(N__45872),
            .in1(N__45462),
            .in2(N__42421),
            .in3(N__45123),
            .lcout(elapsed_time_ns_1_RNI6IU8E1_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_16_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_16_16_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7JU8E1_24_LC_16_16_3  (
            .in0(N__45461),
            .in1(N__45148),
            .in2(N__42436),
            .in3(N__45873),
            .lcout(elapsed_time_ns_1_RNI7JU8E1_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_16_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_16_16_4 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHKEE1_5_LC_16_16_4  (
            .in0(N__42306),
            .in1(N__45460),
            .in2(N__45906),
            .in3(N__42327),
            .lcout(elapsed_time_ns_1_RNIMHKEE1_0_5),
            .ltout(elapsed_time_ns_1_RNIMHKEE1_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_16_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_16_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_16_16_5 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_16_16_5  (
            .in0(N__47076),
            .in1(N__42286),
            .in2(N__42223),
            .in3(N__42216),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49911),
            .ce(N__48951),
            .sr(N__49458));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_16_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_16_16_6 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5IV8E1_31_LC_16_16_6  (
            .in0(N__42136),
            .in1(N__47077),
            .in2(N__45907),
            .in3(N__45464),
            .lcout(elapsed_time_ns_1_RNI5IV8E1_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_16_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_16_17_0 .LUT_INIT=16'b1111110011111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBC0221_19_LC_16_17_0  (
            .in0(N__42962),
            .in1(N__42118),
            .in2(N__45353),
            .in3(N__45514),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_16_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_16_17_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIIC6P1_19_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42103),
            .in3(N__46000),
            .lcout(elapsed_time_ns_1_RNIIIC6P1_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_16_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_16_17_2 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9LU8E1_26_LC_16_17_2  (
            .in0(N__45096),
            .in1(N__42496),
            .in2(N__45549),
            .in3(N__45915),
            .lcout(elapsed_time_ns_1_RNI9LU8E1_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_16_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_16_17_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIBNU8E1_28_LC_16_17_3  (
            .in0(N__45513),
            .in1(N__42546),
            .in2(N__45928),
            .in3(N__42487),
            .lcout(elapsed_time_ns_1_RNIBNU8E1_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_16_17_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_16_17_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAMU8E1_27_LC_16_17_4  (
            .in0(N__42526),
            .in1(N__45911),
            .in2(N__42505),
            .in3(N__45512),
            .lcout(elapsed_time_ns_1_RNIAMU8E1_0_27),
            .ltout(elapsed_time_ns_1_RNIAMU8E1_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_16_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_16_17_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_6_15_LC_16_17_5  (
            .in0(N__42495),
            .in1(N__42486),
            .in2(N__42478),
            .in3(N__42471),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_6Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_16_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_16_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_15_LC_16_17_6  (
            .in0(N__42460),
            .in1(N__42450),
            .in2(N__42439),
            .in3(N__42406),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_16_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_16_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_o5_0_15_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__42432),
            .in2(_gnd_net_),
            .in3(N__42417),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_i_o5_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_16_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_16_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIMHD01_11_LC_16_18_0  (
            .in0(N__45006),
            .in1(N__42399),
            .in2(N__42592),
            .in3(N__42378),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_16_18_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_16_18_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI76C4N_0_31_LC_16_18_1  (
            .in0(N__42367),
            .in1(N__49585),
            .in2(_gnd_net_),
            .in3(N__45313),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_344_i ),
            .ltout(\delay_measurement_inst.delay_hc_timer.N_344_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_16_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_16_18_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIHHC6P1_18_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42352),
            .in3(N__42598),
            .lcout(elapsed_time_ns_1_RNIHHC6P1_0_18),
            .ltout(elapsed_time_ns_1_RNIHHC6P1_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_16_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_16_18_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2_9_LC_16_18_3  (
            .in0(N__42955),
            .in1(N__42773),
            .in2(N__42349),
            .in3(N__42643),
            .lcout(\phase_controller_inst1.stoper_hc.target_time_4_f0_i_o2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_18_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_18_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_16_18_4  (
            .in0(N__42789),
            .in1(N__45801),
            .in2(N__42610),
            .in3(N__42573),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_16_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_16_18_5 .LUT_INIT=16'b1111111010111010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAB0221_18_LC_16_18_5  (
            .in0(N__45315),
            .in1(N__45524),
            .in2(N__43376),
            .in3(N__42609),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_16_18_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_16_18_6 .LUT_INIT=16'b1110111111101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI670221_14_LC_16_18_6  (
            .in0(N__42591),
            .in1(N__45316),
            .in2(N__45550),
            .in3(N__46884),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_16_18_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_16_18_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDDC6P1_14_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42580),
            .in3(N__46013),
            .lcout(elapsed_time_ns_1_RNIDDC6P1_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_16_19_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_16_19_0 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI890221_16_LC_16_19_0  (
            .in0(N__42644),
            .in1(N__45545),
            .in2(N__45352),
            .in3(N__42577),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_16_19_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_16_19_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIFFC6P1_16_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42562),
            .in3(N__46004),
            .lcout(elapsed_time_ns_1_RNIFFC6P1_0_16),
            .ltout(elapsed_time_ns_1_RNIFFC6P1_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_16_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_16_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_16_19_2 .LUT_INIT=16'b0000000011111100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__46794),
            .in2(N__42559),
            .in3(N__47055),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49897),
            .ce(N__49108),
            .sr(N__49482));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_19_3 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_16_19_3  (
            .in0(N__42555),
            .in1(N__48495),
            .in2(N__48523),
            .in3(N__42801),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_19_4 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_19_4  (
            .in0(N__48496),
            .in1(N__48519),
            .in2(N__42805),
            .in3(N__42556),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_16_19_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_16_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_16_19_5 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_16_19_5  (
            .in0(N__47056),
            .in1(_gnd_net_),
            .in2(N__46827),
            .in3(N__42774),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49897),
            .ce(N__49108),
            .sr(N__49482));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_16_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_16_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_16_19_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_16_19_6  (
            .in0(N__42964),
            .in1(N__47057),
            .in2(_gnd_net_),
            .in3(N__46795),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49897),
            .ce(N__49108),
            .sr(N__49482));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_16_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_16_19_7 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_16_19_7  (
            .in0(N__42928),
            .in1(N__48665),
            .in2(N__48475),
            .in3(N__42909),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_16_20_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_16_20_0 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9A0221_17_LC_16_20_0  (
            .in0(N__42769),
            .in1(N__45546),
            .in2(N__45364),
            .in3(N__42793),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_16_20_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_16_20_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIGGC6P1_17_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42778),
            .in3(N__46016),
            .lcout(elapsed_time_ns_1_RNIGGC6P1_0_17),
            .ltout(elapsed_time_ns_1_RNIGGC6P1_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_16_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_16_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_16_20_2 .LUT_INIT=16'b0101010101010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_16_20_2  (
            .in0(N__47059),
            .in1(_gnd_net_),
            .in2(N__42742),
            .in3(N__46810),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49891),
            .ce(N__43148),
            .sr(N__49489));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_16_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_16_20_3 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_16_20_3  (
            .in0(N__42681),
            .in1(N__42618),
            .in2(N__42721),
            .in3(N__42690),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_20_4 .LUT_INIT=16'b0010000011110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_16_20_4  (
            .in0(N__42619),
            .in1(N__42717),
            .in2(N__42694),
            .in3(N__42682),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_16_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_16_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_16_20_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_16_20_5  (
            .in0(N__42645),
            .in1(N__47058),
            .in2(_gnd_net_),
            .in3(N__46799),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49891),
            .ce(N__43148),
            .sr(N__49489));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_16_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_16_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_16_20_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_16_20_6  (
            .in0(N__47060),
            .in1(N__46811),
            .in2(_gnd_net_),
            .in3(N__42963),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49891),
            .ce(N__43148),
            .sr(N__49489));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_16_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_16_21_1 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_i_a2_10_LC_16_21_1  (
            .in0(N__45735),
            .in1(N__46885),
            .in2(_gnd_net_),
            .in3(N__45673),
            .lcout(\phase_controller_inst1.stoper_hc.N_318 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_318_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_16_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_16_21_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_16_21_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_16_21_2  (
            .in0(N__47062),
            .in1(N__43308),
            .in2(N__42931),
            .in3(N__46806),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49883),
            .ce(N__49123),
            .sr(N__49494));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_16_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_16_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_16_21_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_16_21_3  (
            .in0(N__46802),
            .in1(N__47063),
            .in2(N__43264),
            .in3(N__46922),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49883),
            .ce(N__49123),
            .sr(N__49494));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_16_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_16_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_16_21_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_16_21_4  (
            .in0(N__47064),
            .in1(N__46805),
            .in2(N__46930),
            .in3(N__43215),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49883),
            .ce(N__49123),
            .sr(N__49494));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_16_21_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_16_21_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_16_21_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_16_21_5  (
            .in0(N__46803),
            .in1(N__47065),
            .in2(N__44995),
            .in3(N__46923),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49883),
            .ce(N__49123),
            .sr(N__49494));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_16_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_16_21_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_16_21_6 .LUT_INIT=16'b0101010001010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_16_21_6  (
            .in0(N__47061),
            .in1(N__46804),
            .in2(N__43381),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49883),
            .ce(N__49123),
            .sr(N__49494));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_21_7 .LUT_INIT=16'b0100111100000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_21_7  (
            .in0(N__48474),
            .in1(N__42927),
            .in2(N__48673),
            .in3(N__42913),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_22_0 .LUT_INIT=16'b0010001010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_22_0  (
            .in0(N__42894),
            .in1(N__42874),
            .in2(N__43344),
            .in3(N__42850),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_16_22_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_16_22_1 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_16_22_1  (
            .in0(N__47066),
            .in1(N__46822),
            .in2(_gnd_net_),
            .in3(N__43377),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(N__43149),
            .sr(N__49504));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_16_22_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_16_22_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_16_22_2 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_16_22_2  (
            .in0(N__46926),
            .in1(N__47072),
            .in2(N__46831),
            .in3(N__46890),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(N__43149),
            .sr(N__49504));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_16_22_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_16_22_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_16_22_3  (
            .in0(N__47068),
            .in1(N__46927),
            .in2(N__43309),
            .in3(N__46825),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(N__43149),
            .sr(N__49504));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_16_22_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_16_22_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_16_22_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_16_22_4  (
            .in0(N__46924),
            .in1(N__47069),
            .in2(N__46829),
            .in3(N__43263),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(N__43149),
            .sr(N__49504));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_16_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_16_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_16_22_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_16_22_5  (
            .in0(N__47070),
            .in1(N__46823),
            .in2(N__43219),
            .in3(N__46928),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(N__43149),
            .sr(N__49504));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_16_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_16_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_16_22_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_16_22_6  (
            .in0(N__46925),
            .in1(N__47071),
            .in2(N__46830),
            .in3(N__44994),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(N__43149),
            .sr(N__49504));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_16_22_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_16_22_7 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_16_22_7  (
            .in0(N__47067),
            .in1(N__45756),
            .in2(N__45610),
            .in3(N__46824),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49877),
            .ce(N__43149),
            .sr(N__49504));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_17_7_0  (
            .in0(N__43822),
            .in1(N__46520),
            .in2(_gnd_net_),
            .in3(N__42970),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__49966),
            .ce(N__43687),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_17_7_1  (
            .in0(N__43818),
            .in1(N__47498),
            .in2(_gnd_net_),
            .in3(N__42967),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__49966),
            .ce(N__43687),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_17_7_2  (
            .in0(N__43823),
            .in1(N__43620),
            .in2(_gnd_net_),
            .in3(N__43408),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__49966),
            .ce(N__43687),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_17_7_3  (
            .in0(N__43819),
            .in1(N__43596),
            .in2(_gnd_net_),
            .in3(N__43405),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__49966),
            .ce(N__43687),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_17_7_4  (
            .in0(N__43824),
            .in1(N__43571),
            .in2(_gnd_net_),
            .in3(N__43402),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__49966),
            .ce(N__43687),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_17_7_5  (
            .in0(N__43820),
            .in1(N__43544),
            .in2(_gnd_net_),
            .in3(N__43399),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__49966),
            .ce(N__43687),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_17_7_6  (
            .in0(N__43825),
            .in1(N__43518),
            .in2(_gnd_net_),
            .in3(N__43396),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__49966),
            .ce(N__43687),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_17_7_7  (
            .in0(N__43821),
            .in1(N__43494),
            .in2(_gnd_net_),
            .in3(N__43393),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__49966),
            .ce(N__43687),
            .sr(N__49407));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_17_8_0  (
            .in0(N__43772),
            .in1(N__44120),
            .in2(_gnd_net_),
            .in3(N__43390),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__49961),
            .ce(N__43683),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_17_8_1  (
            .in0(N__43776),
            .in1(N__44072),
            .in2(_gnd_net_),
            .in3(N__43387),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__49961),
            .ce(N__43683),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_17_8_2  (
            .in0(N__43769),
            .in1(N__44025),
            .in2(_gnd_net_),
            .in3(N__43384),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__49961),
            .ce(N__43683),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_17_8_3  (
            .in0(N__43773),
            .in1(N__43973),
            .in2(_gnd_net_),
            .in3(N__43435),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__49961),
            .ce(N__43683),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_17_8_4  (
            .in0(N__43770),
            .in1(N__43946),
            .in2(_gnd_net_),
            .in3(N__43432),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__49961),
            .ce(N__43683),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_17_8_5  (
            .in0(N__43774),
            .in1(N__43898),
            .in2(_gnd_net_),
            .in3(N__43429),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__49961),
            .ce(N__43683),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_17_8_6  (
            .in0(N__43771),
            .in1(N__43872),
            .in2(_gnd_net_),
            .in3(N__43426),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__49961),
            .ce(N__43683),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_17_8_7  (
            .in0(N__43775),
            .in1(N__43842),
            .in2(_gnd_net_),
            .in3(N__43423),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__49961),
            .ce(N__43683),
            .sr(N__49409));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_17_9_0  (
            .in0(N__43777),
            .in1(N__44462),
            .in2(_gnd_net_),
            .in3(N__43420),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__49955),
            .ce(N__43676),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_17_9_1  (
            .in0(N__43814),
            .in1(N__44435),
            .in2(_gnd_net_),
            .in3(N__43417),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__49955),
            .ce(N__43676),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_17_9_2  (
            .in0(N__43778),
            .in1(N__44393),
            .in2(_gnd_net_),
            .in3(N__43414),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__49955),
            .ce(N__43676),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_17_9_3  (
            .in0(N__43815),
            .in1(N__44354),
            .in2(_gnd_net_),
            .in3(N__43411),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__49955),
            .ce(N__43676),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_17_9_4  (
            .in0(N__43779),
            .in1(N__44309),
            .in2(_gnd_net_),
            .in3(N__43462),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__49955),
            .ce(N__43676),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_17_9_5  (
            .in0(N__43816),
            .in1(N__44264),
            .in2(_gnd_net_),
            .in3(N__43459),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__49955),
            .ce(N__43676),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_17_9_6  (
            .in0(N__43780),
            .in1(N__44220),
            .in2(_gnd_net_),
            .in3(N__43456),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__49955),
            .ce(N__43676),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_17_9_7  (
            .in0(N__43817),
            .in1(N__44175),
            .in2(_gnd_net_),
            .in3(N__43453),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__49955),
            .ce(N__43676),
            .sr(N__49411));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_17_10_0  (
            .in0(N__43808),
            .in1(N__44933),
            .in2(_gnd_net_),
            .in3(N__43450),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__49950),
            .ce(N__43675),
            .sr(N__49413));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_17_10_1  (
            .in0(N__43812),
            .in1(N__44876),
            .in2(_gnd_net_),
            .in3(N__43447),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__49950),
            .ce(N__43675),
            .sr(N__49413));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_17_10_2  (
            .in0(N__43809),
            .in1(N__44804),
            .in2(_gnd_net_),
            .in3(N__43444),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__49950),
            .ce(N__43675),
            .sr(N__49413));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_17_10_3  (
            .in0(N__43813),
            .in1(N__44758),
            .in2(_gnd_net_),
            .in3(N__43441),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__49950),
            .ce(N__43675),
            .sr(N__49413));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_17_10_4  (
            .in0(N__43810),
            .in1(N__44823),
            .in2(_gnd_net_),
            .in3(N__43438),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__49950),
            .ce(N__43675),
            .sr(N__49413));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_17_10_5  (
            .in0(N__44736),
            .in1(N__43811),
            .in2(_gnd_net_),
            .in3(N__43690),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49950),
            .ce(N__43675),
            .sr(N__49413));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__43626),
            .in2(N__46534),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__49946),
            .ce(N__47475),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__43602),
            .in2(N__47512),
            .in3(N__43630),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__49946),
            .ce(N__47475),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__43627),
            .in2(N__43578),
            .in3(N__43606),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__49946),
            .ce(N__47475),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__43603),
            .in2(N__43551),
            .in3(N__43582),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__49946),
            .ce(N__47475),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__43524),
            .in2(N__43579),
            .in3(N__43555),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__49946),
            .ce(N__47475),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__43500),
            .in2(N__43552),
            .in3(N__43528),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__49946),
            .ce(N__47475),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__43525),
            .in2(N__44127),
            .in3(N__43504),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__49946),
            .ce(N__47475),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__43501),
            .in2(N__44079),
            .in3(N__43465),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__49946),
            .ce(N__47475),
            .sr(N__49416));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__44031),
            .in2(N__44131),
            .in3(N__44083),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__49941),
            .ce(N__47477),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__43980),
            .in2(N__44080),
            .in3(N__44035),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__49941),
            .ce(N__47477),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__44032),
            .in2(N__43953),
            .in3(N__43990),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__49941),
            .ce(N__47477),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__43899),
            .in2(N__43987),
            .in3(N__43957),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__49941),
            .ce(N__47477),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__43878),
            .in2(N__43954),
            .in3(N__43903),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr9lto15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__49941),
            .ce(N__47477),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(N__43900),
            .in2(N__43854),
            .in3(N__43882),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__49941),
            .ce(N__47477),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__43879),
            .in2(N__44475),
            .in3(N__43858),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__49941),
            .ce(N__47477),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__44436),
            .in2(N__43855),
            .in3(N__43828),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__49941),
            .ce(N__47477),
            .sr(N__49423));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__44394),
            .in2(N__44476),
            .in3(N__44446),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__49934),
            .ce(N__47478),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__44355),
            .in2(N__44443),
            .in3(N__44398),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__49934),
            .ce(N__47478),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__44395),
            .in2(N__44316),
            .in3(N__44359),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__49934),
            .ce(N__47478),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__44356),
            .in2(N__44271),
            .in3(N__44320),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__49934),
            .ce(N__47478),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(N__44226),
            .in2(N__44317),
            .in3(N__44275),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__49934),
            .ce(N__47478),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__44181),
            .in2(N__44272),
            .in3(N__44230),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__49934),
            .ce(N__47478),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(N__44227),
            .in2(N__44940),
            .in3(N__44185),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__49934),
            .ce(N__47478),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_17_13_7  (
            .in0(_gnd_net_),
            .in1(N__44182),
            .in2(N__44883),
            .in3(N__44134),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__49934),
            .ce(N__47478),
            .sr(N__49425));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__44805),
            .in2(N__44941),
            .in3(N__44890),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__49929),
            .ce(N__47479),
            .sr(N__49435));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__44756),
            .in2(N__44887),
            .in3(N__44827),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__49929),
            .ce(N__47479),
            .sr(N__49435));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__44824),
            .in2(N__44809),
            .in3(N__44761),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__49929),
            .ce(N__47479),
            .sr(N__49435));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(N__44757),
            .in2(N__44740),
            .in3(N__44701),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__49929),
            .ce(N__47479),
            .sr(N__49435));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44698),
            .lcout(\delay_measurement_inst.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49929),
            .ce(N__47479),
            .sr(N__49435));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_17_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_17_15_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_17_15_0  (
            .in0(N__44641),
            .in1(N__46665),
            .in2(N__46606),
            .in3(N__44597),
            .lcout(),
            .ltout(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_LC_17_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_17_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_17_15_1 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_17_15_1  (
            .in0(N__44557),
            .in1(N__44503),
            .in2(N__44479),
            .in3(N__50131),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49923),
            .ce(),
            .sr(N__49441));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_17_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_17_15_4 .LUT_INIT=16'b1111011111110101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNID27N1_28_LC_17_15_4  (
            .in0(N__50106),
            .in1(N__48200),
            .in2(N__48171),
            .in3(N__45196),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_15_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45187),
            .in3(N__50017),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_17_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_17_15_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2_28_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__50018),
            .in2(_gnd_net_),
            .in3(N__45180),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIJF7V2Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_17_16_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_17_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI22I01_23_LC_17_16_0  (
            .in0(N__45168),
            .in1(N__45147),
            .in2(N__45127),
            .in3(N__45097),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_17_16_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_17_16_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPFU14_11_LC_17_16_1  (
            .in0(N__45076),
            .in1(N__45070),
            .in2(N__45058),
            .in3(N__45055),
            .lcout(\delay_measurement_inst.delay_hc_timer.un6_elapsed_time_trlto30_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_16_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_17_16_2  (
            .in0(N__48231),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48216),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_16_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_17_16_3  (
            .in0(N__48261),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48246),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_17_16_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_17_16_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI5GT8E1_13_LC_17_16_4  (
            .in0(N__45013),
            .in1(N__45922),
            .in2(N__44987),
            .in3(N__45470),
            .lcout(elapsed_time_ns_1_RNI5GT8E1_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_17_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_17_16_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_17_16_5  (
            .in0(_gnd_net_),
            .in1(N__48166),
            .in2(_gnd_net_),
            .in3(N__48201),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_17_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_17_17_0 .LUT_INIT=16'b1111111010101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIN8N721_6_LC_17_17_0  (
            .in0(N__45374),
            .in1(N__45958),
            .in2(N__45552),
            .in3(N__46047),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_17_17_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_17_17_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUE3CP1_6_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46027),
            .in3(N__46014),
            .lcout(elapsed_time_ns_1_RNIUE3CP1_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_17_17_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_17_17_2 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7IT8E1_15_LC_17_17_2  (
            .in0(N__45701),
            .in1(N__45926),
            .in2(N__45551),
            .in3(N__45808),
            .lcout(elapsed_time_ns_1_RNI7IT8E1_0_15),
            .ltout(elapsed_time_ns_1_RNI7IT8E1_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.N_269_i_1_LC_17_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.N_269_i_1_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.N_269_i_1_LC_17_17_3 .LUT_INIT=16'b0101000001010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.N_269_i_1_LC_17_17_3  (
            .in0(N__45654),
            .in1(N__46870),
            .in2(N__45790),
            .in3(N__45779),
            .lcout(\phase_controller_inst1.stoper_hc.N_269_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_17_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_17_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_17_17_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_17_17_6  (
            .in0(N__47020),
            .in1(N__46745),
            .in2(N__45717),
            .in3(N__45655),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49912),
            .ce(N__48993),
            .sr(N__49459));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_17_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_17_17_7 .LUT_INIT=16'b1111111110101100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQBN721_9_LC_17_17_7  (
            .in0(N__45630),
            .in1(N__45609),
            .in2(N__45556),
            .in3(N__45375),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc_1_latch_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_17_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_17_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__46218),
            .in2(_gnd_net_),
            .in3(N__46245),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_17_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_17_18_1 .LUT_INIT=16'b1111011111110101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI5B3T_28_LC_17_18_1  (
            .in0(N__46126),
            .in1(N__48736),
            .in2(N__48715),
            .in3(N__47140),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_17_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_17_18_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1_28_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46252),
            .in3(N__46219),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNITOIN1Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_17_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_17_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_17_18_3 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_17_18_3  (
            .in0(N__46220),
            .in1(N__48994),
            .in2(N__46249),
            .in3(N__48142),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49907),
            .ce(),
            .sr(N__49465));
    defparam \phase_controller_inst2.stoper_hc.running_LC_17_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_17_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_17_18_4 .LUT_INIT=16'b1011001111110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_17_18_4  (
            .in0(N__47124),
            .in1(N__46127),
            .in2(N__46237),
            .in3(N__46221),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49907),
            .ce(),
            .sr(N__49465));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_17_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_17_18_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_17_18_5  (
            .in0(N__46125),
            .in1(N__46233),
            .in2(_gnd_net_),
            .in3(N__46158),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_17_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_17_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_17_18_6 .LUT_INIT=16'b1101110000001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_17_18_6  (
            .in0(N__47125),
            .in1(N__46181),
            .in2(N__46225),
            .in3(N__46128),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49907),
            .ce(),
            .sr(N__49465));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_17_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_17_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_17_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46159),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49907),
            .ce(),
            .sr(N__49465));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_17_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_17_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__46108),
            .in2(N__46099),
            .in3(N__48140),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_17_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_17_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__46090),
            .in2(N__46078),
            .in3(N__48115),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_17_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_17_19_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_17_19_2  (
            .in0(N__48435),
            .in1(N__46069),
            .in2(N__46057),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_17_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_17_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__46411),
            .in2(N__46402),
            .in3(N__48415),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_17_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_17_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__46393),
            .in2(N__46381),
            .in3(N__48397),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_17_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_17_19_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_17_19_5  (
            .in0(N__48379),
            .in1(N__46369),
            .in2(N__46354),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_17_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_17_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__46345),
            .in2(N__46330),
            .in3(N__48361),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_17_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_17_19_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_17_19_7  (
            .in0(N__48343),
            .in1(N__46318),
            .in2(N__46309),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_17_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_17_20_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_17_20_0  (
            .in0(N__48325),
            .in1(N__46300),
            .in2(N__46291),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_17_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_17_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__46282),
            .in2(N__46276),
            .in3(N__48307),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_17_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_17_20_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_17_20_2  (
            .in0(N__48616),
            .in1(N__46267),
            .in2(N__46261),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_17_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_17_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__46492),
            .in2(N__46501),
            .in3(N__48595),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_17_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_17_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__46486),
            .in2(N__46480),
            .in3(N__48577),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_17_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_17_20_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_17_20_5  (
            .in0(N__48559),
            .in1(N__46471),
            .in2(N__46678),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_17_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_17_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__46465),
            .in2(N__46456),
            .in3(N__48541),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_17_20_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_17_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(N__46447),
            .in2(N__46441),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_17_21_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_17_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(N__46429),
            .in2(N__46420),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_17_21_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_17_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(N__50329),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_17_21_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_17_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__48772),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_17_21_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_17_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(N__50365),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_17_21_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_17_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(N__48808),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_17_21_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_17_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(N__48742),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_21_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(N__48679),
            .in2(N__48711),
            .in3(N__47131),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47128),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_17_22_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_17_22_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_17_22_5 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_17_22_5  (
            .in0(N__47113),
            .in1(N__46929),
            .in2(N__46891),
            .in3(N__46828),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49884),
            .ce(N__49069),
            .sr(N__49495));
    defparam \phase_controller_inst1.T12_LC_17_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.T12_LC_17_23_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T12_LC_17_23_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst1.T12_LC_17_23_1  (
            .in0(N__46545),
            .in1(N__46666),
            .in2(_gnd_net_),
            .in3(N__46599),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49878),
            .ce(),
            .sr(N__49505));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46533),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(N__47476),
            .sr(N__49412));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47511),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49956),
            .ce(N__47476),
            .sr(N__49412));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_18_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_18_11_0 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNINAPP_2_LC_18_11_0  (
            .in0(N__47382),
            .in1(N__47762),
            .in2(N__47364),
            .in3(N__47791),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_19_LC_18_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_19_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_19_LC_18_11_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIBHFU2_19_LC_18_11_1  (
            .in0(N__47172),
            .in1(N__47428),
            .in2(N__47458),
            .in3(N__47395),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2BNE1_16_LC_18_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2BNE1_16_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2BNE1_16_LC_18_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2BNE1_16_LC_18_11_2  (
            .in0(N__47226),
            .in1(N__47189),
            .in2(N__47742),
            .in3(N__47207),
            .lcout(\delay_measurement_inst.delay_tr_timer.un1_delay_tr_0_sqmuxa_i_a2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_18_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_18_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJ7L7_4_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(N__47421),
            .in2(_gnd_net_),
            .in3(N__47406),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_346 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_18_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_18_11_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI8R4J_1_LC_18_11_4  (
            .in0(N__47381),
            .in1(N__47351),
            .in2(N__47335),
            .in3(N__47322),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_349 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_349_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_18_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_18_11_5 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_18_11_5  (
            .in0(N__47291),
            .in1(N__47264),
            .in2(N__47248),
            .in3(N__47734),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_11_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIM96P1_16_LC_18_11_6  (
            .in0(N__47225),
            .in1(N__47208),
            .in2(N__47194),
            .in3(N__47171),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_362 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.N_362_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_18_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_18_11_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI965F2_6_LC_18_11_7  (
            .in0(N__47792),
            .in1(N__47763),
            .in2(N__47746),
            .in3(N__47738),
            .lcout(\delay_measurement_inst.N_365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__47689),
            .in2(N__47680),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_18_13_1  (
            .in0(N__50288),
            .in1(N__47655),
            .in2(_gnd_net_),
            .in3(N__47641),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_13_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_18_13_2  (
            .in0(N__50293),
            .in1(N__47622),
            .in2(N__47638),
            .in3(N__47608),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_18_13_3  (
            .in0(N__50289),
            .in1(N__47601),
            .in2(_gnd_net_),
            .in3(N__47587),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_18_13_4  (
            .in0(N__50294),
            .in1(N__47583),
            .in2(_gnd_net_),
            .in3(N__47569),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_18_13_5  (
            .in0(N__50290),
            .in1(N__47565),
            .in2(_gnd_net_),
            .in3(N__47551),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_18_13_6  (
            .in0(N__50295),
            .in1(N__47544),
            .in2(_gnd_net_),
            .in3(N__47530),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_18_13_7  (
            .in0(N__50291),
            .in1(N__47526),
            .in2(_gnd_net_),
            .in3(N__47944),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__49942),
            .ce(),
            .sr(N__49424));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_18_14_0  (
            .in0(N__50276),
            .in1(N__47940),
            .in2(_gnd_net_),
            .in3(N__47926),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_18_14_1  (
            .in0(N__50269),
            .in1(N__47922),
            .in2(_gnd_net_),
            .in3(N__47908),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_18_14_2  (
            .in0(N__50273),
            .in1(N__47904),
            .in2(_gnd_net_),
            .in3(N__47890),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_18_14_3  (
            .in0(N__50270),
            .in1(N__47886),
            .in2(_gnd_net_),
            .in3(N__47872),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_18_14_4  (
            .in0(N__50274),
            .in1(N__47868),
            .in2(_gnd_net_),
            .in3(N__47854),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_18_14_5  (
            .in0(N__50271),
            .in1(N__47850),
            .in2(_gnd_net_),
            .in3(N__47836),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_18_14_6  (
            .in0(N__50275),
            .in1(N__47832),
            .in2(_gnd_net_),
            .in3(N__47818),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_18_14_7  (
            .in0(N__50272),
            .in1(N__47813),
            .in2(_gnd_net_),
            .in3(N__47797),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__49935),
            .ce(),
            .sr(N__49426));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_18_15_0  (
            .in0(N__50277),
            .in1(N__48087),
            .in2(_gnd_net_),
            .in3(N__48073),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__49930),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_18_15_1  (
            .in0(N__50281),
            .in1(N__48063),
            .in2(_gnd_net_),
            .in3(N__48049),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__49930),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_18_15_2  (
            .in0(N__50278),
            .in1(N__48036),
            .in2(_gnd_net_),
            .in3(N__48022),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__49930),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_18_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_18_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_18_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_18_15_3  (
            .in0(N__50282),
            .in1(N__48861),
            .in2(_gnd_net_),
            .in3(N__48019),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__49930),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_18_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_18_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_18_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_18_15_4  (
            .in0(N__50279),
            .in1(N__48876),
            .in2(_gnd_net_),
            .in3(N__48016),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__49930),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_18_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_18_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_18_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_18_15_5  (
            .in0(N__50283),
            .in1(N__48009),
            .in2(_gnd_net_),
            .in3(N__47995),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__49930),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_18_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_18_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_18_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_18_15_6  (
            .in0(N__50280),
            .in1(N__47985),
            .in2(_gnd_net_),
            .in3(N__47971),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__49930),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_18_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_18_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_18_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_18_15_7  (
            .in0(N__50284),
            .in1(N__47961),
            .in2(_gnd_net_),
            .in3(N__47947),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__49930),
            .ce(),
            .sr(N__49436));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_18_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_18_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_18_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_18_16_0  (
            .in0(N__50301),
            .in1(N__48279),
            .in2(_gnd_net_),
            .in3(N__48265),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49442));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_18_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_18_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_18_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_18_16_1  (
            .in0(N__50305),
            .in1(N__48262),
            .in2(_gnd_net_),
            .in3(N__48250),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49442));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_18_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_18_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_18_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_18_16_2  (
            .in0(N__50302),
            .in1(N__48247),
            .in2(_gnd_net_),
            .in3(N__48235),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49442));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_18_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_18_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_18_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_18_16_3  (
            .in0(N__50306),
            .in1(N__48232),
            .in2(_gnd_net_),
            .in3(N__48220),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49442));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_18_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_18_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_18_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_18_16_4  (
            .in0(N__50303),
            .in1(N__48217),
            .in2(_gnd_net_),
            .in3(N__48205),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49442));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_18_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_18_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_18_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_18_16_5  (
            .in0(N__50307),
            .in1(N__48202),
            .in2(_gnd_net_),
            .in3(N__48184),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__49924),
            .ce(),
            .sr(N__49442));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_18_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_18_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_18_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_18_16_6  (
            .in0(N__50304),
            .in1(N__48170),
            .in2(_gnd_net_),
            .in3(N__48181),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49924),
            .ce(),
            .sr(N__49442));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__48141),
            .in2(N__48124),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_18_17_1  (
            .in0(N__48983),
            .in1(N__48114),
            .in2(_gnd_net_),
            .in3(N__48100),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_17_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_18_17_2  (
            .in0(N__48961),
            .in1(N__48442),
            .in2(N__48436),
            .in3(N__48418),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_18_17_3  (
            .in0(N__48984),
            .in1(N__48414),
            .in2(_gnd_net_),
            .in3(N__48400),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_18_17_4  (
            .in0(N__48962),
            .in1(N__48396),
            .in2(_gnd_net_),
            .in3(N__48382),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_18_17_5  (
            .in0(N__48985),
            .in1(N__48378),
            .in2(_gnd_net_),
            .in3(N__48364),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_18_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_18_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_18_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_18_17_6  (
            .in0(N__48963),
            .in1(N__48360),
            .in2(_gnd_net_),
            .in3(N__48346),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_18_17_7  (
            .in0(N__48986),
            .in1(N__48342),
            .in2(_gnd_net_),
            .in3(N__48328),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__49917),
            .ce(),
            .sr(N__49451));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_18_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_18_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_18_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_18_18_0  (
            .in0(N__49104),
            .in1(N__48324),
            .in2(_gnd_net_),
            .in3(N__48310),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__49913),
            .ce(),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_18_18_1  (
            .in0(N__49079),
            .in1(N__48303),
            .in2(_gnd_net_),
            .in3(N__48289),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__49913),
            .ce(),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_18_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_18_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_18_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_18_18_2  (
            .in0(N__49101),
            .in1(N__48615),
            .in2(_gnd_net_),
            .in3(N__48598),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__49913),
            .ce(),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_18_18_3  (
            .in0(N__49080),
            .in1(N__48594),
            .in2(_gnd_net_),
            .in3(N__48580),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__49913),
            .ce(),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_18_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_18_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_18_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_18_18_4  (
            .in0(N__49102),
            .in1(N__48576),
            .in2(_gnd_net_),
            .in3(N__48562),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__49913),
            .ce(),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_18_18_5  (
            .in0(N__49081),
            .in1(N__48558),
            .in2(_gnd_net_),
            .in3(N__48544),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__49913),
            .ce(),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_18_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_18_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_18_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_18_18_6  (
            .in0(N__49103),
            .in1(N__48540),
            .in2(_gnd_net_),
            .in3(N__48526),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__49913),
            .ce(),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_18_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_18_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_18_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_18_18_7  (
            .in0(N__49082),
            .in1(N__48513),
            .in2(_gnd_net_),
            .in3(N__48499),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__49913),
            .ce(),
            .sr(N__49460));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_18_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_18_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_18_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_18_19_0  (
            .in0(N__49083),
            .in1(N__48494),
            .in2(_gnd_net_),
            .in3(N__48478),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__49908),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_18_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_18_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_18_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_18_19_1  (
            .in0(N__49087),
            .in1(N__48467),
            .in2(_gnd_net_),
            .in3(N__48445),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__49908),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_18_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_18_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_18_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_18_19_2  (
            .in0(N__49084),
            .in1(N__48669),
            .in2(_gnd_net_),
            .in3(N__48643),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__49908),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_18_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_18_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_18_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_18_19_3  (
            .in0(N__49088),
            .in1(N__50343),
            .in2(_gnd_net_),
            .in3(N__48640),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__49908),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_18_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_18_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_18_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_18_19_4  (
            .in0(N__49085),
            .in1(N__50358),
            .in2(_gnd_net_),
            .in3(N__48637),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__49908),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_18_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_18_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_18_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_18_19_5  (
            .in0(N__49089),
            .in1(N__48786),
            .in2(_gnd_net_),
            .in3(N__48634),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__49908),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_18_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_18_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_18_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_18_19_6  (
            .in0(N__49086),
            .in1(N__48801),
            .in2(_gnd_net_),
            .in3(N__48631),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__49908),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_18_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_18_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_18_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_18_19_7  (
            .in0(N__49090),
            .in1(N__50379),
            .in2(_gnd_net_),
            .in3(N__48628),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__49908),
            .ce(),
            .sr(N__49466));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_18_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_18_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_18_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_18_20_0  (
            .in0(N__49098),
            .in1(N__50392),
            .in2(_gnd_net_),
            .in3(N__48625),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__49902),
            .ce(),
            .sr(N__49473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_18_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_18_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_18_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_18_20_1  (
            .in0(N__49091),
            .in1(N__48820),
            .in2(_gnd_net_),
            .in3(N__48622),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__49902),
            .ce(),
            .sr(N__49473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_18_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_18_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_18_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_18_20_2  (
            .in0(N__49099),
            .in1(N__48832),
            .in2(_gnd_net_),
            .in3(N__48619),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__49902),
            .ce(),
            .sr(N__49473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_18_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_18_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_18_20_3  (
            .in0(N__49092),
            .in1(N__48754),
            .in2(_gnd_net_),
            .in3(N__49132),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__49902),
            .ce(),
            .sr(N__49473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_18_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_18_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_18_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_18_20_4  (
            .in0(N__49100),
            .in1(N__48766),
            .in2(_gnd_net_),
            .in3(N__49129),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__49902),
            .ce(),
            .sr(N__49473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_18_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_18_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_18_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_18_20_5  (
            .in0(N__49093),
            .in1(N__48735),
            .in2(_gnd_net_),
            .in3(N__49126),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__49902),
            .ce(),
            .sr(N__49473));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_18_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_18_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_18_20_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_18_20_6  (
            .in0(N__48706),
            .in1(N__49094),
            .in2(_gnd_net_),
            .in3(N__48883),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49902),
            .ce(),
            .sr(N__49473));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_18_21_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_18_21_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__48880),
            .in2(_gnd_net_),
            .in3(N__48862),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_21_1  (
            .in0(_gnd_net_),
            .in1(N__48831),
            .in2(_gnd_net_),
            .in3(N__48819),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_18_21_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_18_21_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(N__48802),
            .in2(_gnd_net_),
            .in3(N__48787),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_21_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_18_21_3  (
            .in0(_gnd_net_),
            .in1(N__48765),
            .in2(_gnd_net_),
            .in3(N__48753),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_21_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_18_21_4  (
            .in0(N__48734),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48710),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_21_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_21_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_21_6  (
            .in0(_gnd_net_),
            .in1(N__50391),
            .in2(_gnd_net_),
            .in3(N__50380),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_21_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_21_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_21_7  (
            .in0(_gnd_net_),
            .in1(N__50359),
            .in2(_gnd_net_),
            .in3(N__50344),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_df20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_14_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_14_6  (
            .in0(_gnd_net_),
            .in1(N__50102),
            .in2(_gnd_net_),
            .in3(N__50139),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_20_15_5  (
            .in0(N__50088),
            .in1(N__49989),
            .in2(_gnd_net_),
            .in3(N__50132),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_20_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_20_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_20_16_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_20_16_1  (
            .in0(N__50140),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49936),
            .ce(),
            .sr(N__49443));
    defparam \phase_controller_inst1.stoper_tr.running_LC_20_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_20_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_20_16_5 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_20_16_5  (
            .in0(N__50098),
            .in1(N__50062),
            .in2(N__49993),
            .in3(N__50016),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49936),
            .ce(),
            .sr(N__49443));
endmodule // MAIN
