// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 2 2025 23:51:13

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    start_stop,
    s2_phy,
    T23,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    T45,
    T12,
    s4_phy,
    rgb_g,
    T01,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    input start_stop;
    output s2_phy;
    output T23;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output T45;
    output T12;
    output s4_phy;
    output rgb_g;
    output T01;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__48452;
    wire N__48451;
    wire N__48450;
    wire N__48441;
    wire N__48440;
    wire N__48439;
    wire N__48432;
    wire N__48431;
    wire N__48430;
    wire N__48423;
    wire N__48422;
    wire N__48421;
    wire N__48414;
    wire N__48413;
    wire N__48412;
    wire N__48405;
    wire N__48404;
    wire N__48403;
    wire N__48396;
    wire N__48395;
    wire N__48394;
    wire N__48387;
    wire N__48386;
    wire N__48385;
    wire N__48378;
    wire N__48377;
    wire N__48376;
    wire N__48369;
    wire N__48368;
    wire N__48367;
    wire N__48360;
    wire N__48359;
    wire N__48358;
    wire N__48351;
    wire N__48350;
    wire N__48349;
    wire N__48342;
    wire N__48341;
    wire N__48340;
    wire N__48333;
    wire N__48332;
    wire N__48331;
    wire N__48324;
    wire N__48323;
    wire N__48322;
    wire N__48315;
    wire N__48314;
    wire N__48313;
    wire N__48306;
    wire N__48305;
    wire N__48304;
    wire N__48287;
    wire N__48286;
    wire N__48285;
    wire N__48284;
    wire N__48281;
    wire N__48278;
    wire N__48275;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48263;
    wire N__48260;
    wire N__48257;
    wire N__48254;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48242;
    wire N__48239;
    wire N__48236;
    wire N__48227;
    wire N__48226;
    wire N__48223;
    wire N__48222;
    wire N__48219;
    wire N__48216;
    wire N__48213;
    wire N__48206;
    wire N__48205;
    wire N__48204;
    wire N__48203;
    wire N__48202;
    wire N__48201;
    wire N__48200;
    wire N__48199;
    wire N__48198;
    wire N__48197;
    wire N__48196;
    wire N__48195;
    wire N__48194;
    wire N__48193;
    wire N__48190;
    wire N__48189;
    wire N__48188;
    wire N__48187;
    wire N__48186;
    wire N__48185;
    wire N__48184;
    wire N__48183;
    wire N__48182;
    wire N__48181;
    wire N__48180;
    wire N__48179;
    wire N__48178;
    wire N__48177;
    wire N__48176;
    wire N__48173;
    wire N__48170;
    wire N__48169;
    wire N__48160;
    wire N__48155;
    wire N__48154;
    wire N__48153;
    wire N__48152;
    wire N__48151;
    wire N__48150;
    wire N__48149;
    wire N__48148;
    wire N__48147;
    wire N__48146;
    wire N__48145;
    wire N__48144;
    wire N__48133;
    wire N__48132;
    wire N__48131;
    wire N__48130;
    wire N__48129;
    wire N__48118;
    wire N__48117;
    wire N__48116;
    wire N__48105;
    wire N__48102;
    wire N__48101;
    wire N__48100;
    wire N__48099;
    wire N__48098;
    wire N__48097;
    wire N__48096;
    wire N__48095;
    wire N__48092;
    wire N__48091;
    wire N__48090;
    wire N__48089;
    wire N__48088;
    wire N__48087;
    wire N__48080;
    wire N__48073;
    wire N__48068;
    wire N__48063;
    wire N__48060;
    wire N__48057;
    wire N__48052;
    wire N__48051;
    wire N__48042;
    wire N__48039;
    wire N__48036;
    wire N__48027;
    wire N__48026;
    wire N__48025;
    wire N__48024;
    wire N__48023;
    wire N__48022;
    wire N__48021;
    wire N__48020;
    wire N__48019;
    wire N__48016;
    wire N__48011;
    wire N__48010;
    wire N__48009;
    wire N__48008;
    wire N__48007;
    wire N__48006;
    wire N__48005;
    wire N__48004;
    wire N__48003;
    wire N__48002;
    wire N__48001;
    wire N__48000;
    wire N__47999;
    wire N__47998;
    wire N__47997;
    wire N__47996;
    wire N__47995;
    wire N__47992;
    wire N__47989;
    wire N__47988;
    wire N__47987;
    wire N__47986;
    wire N__47985;
    wire N__47984;
    wire N__47983;
    wire N__47982;
    wire N__47981;
    wire N__47980;
    wire N__47971;
    wire N__47960;
    wire N__47951;
    wire N__47936;
    wire N__47933;
    wire N__47928;
    wire N__47925;
    wire N__47922;
    wire N__47917;
    wire N__47910;
    wire N__47903;
    wire N__47898;
    wire N__47895;
    wire N__47886;
    wire N__47879;
    wire N__47870;
    wire N__47861;
    wire N__47856;
    wire N__47853;
    wire N__47848;
    wire N__47839;
    wire N__47834;
    wire N__47827;
    wire N__47824;
    wire N__47813;
    wire N__47806;
    wire N__47777;
    wire N__47776;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47766;
    wire N__47763;
    wire N__47762;
    wire N__47759;
    wire N__47756;
    wire N__47753;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47741;
    wire N__47738;
    wire N__47735;
    wire N__47730;
    wire N__47723;
    wire N__47722;
    wire N__47719;
    wire N__47718;
    wire N__47715;
    wire N__47712;
    wire N__47709;
    wire N__47702;
    wire N__47701;
    wire N__47700;
    wire N__47699;
    wire N__47698;
    wire N__47697;
    wire N__47696;
    wire N__47695;
    wire N__47694;
    wire N__47693;
    wire N__47692;
    wire N__47691;
    wire N__47690;
    wire N__47689;
    wire N__47688;
    wire N__47687;
    wire N__47686;
    wire N__47685;
    wire N__47684;
    wire N__47683;
    wire N__47682;
    wire N__47681;
    wire N__47680;
    wire N__47679;
    wire N__47678;
    wire N__47677;
    wire N__47676;
    wire N__47675;
    wire N__47674;
    wire N__47673;
    wire N__47672;
    wire N__47671;
    wire N__47670;
    wire N__47669;
    wire N__47668;
    wire N__47667;
    wire N__47666;
    wire N__47665;
    wire N__47664;
    wire N__47663;
    wire N__47662;
    wire N__47661;
    wire N__47660;
    wire N__47659;
    wire N__47658;
    wire N__47657;
    wire N__47656;
    wire N__47655;
    wire N__47654;
    wire N__47653;
    wire N__47652;
    wire N__47651;
    wire N__47650;
    wire N__47649;
    wire N__47648;
    wire N__47647;
    wire N__47646;
    wire N__47645;
    wire N__47644;
    wire N__47643;
    wire N__47642;
    wire N__47641;
    wire N__47640;
    wire N__47639;
    wire N__47638;
    wire N__47637;
    wire N__47636;
    wire N__47635;
    wire N__47634;
    wire N__47633;
    wire N__47632;
    wire N__47631;
    wire N__47630;
    wire N__47629;
    wire N__47628;
    wire N__47627;
    wire N__47626;
    wire N__47625;
    wire N__47624;
    wire N__47623;
    wire N__47622;
    wire N__47621;
    wire N__47620;
    wire N__47619;
    wire N__47618;
    wire N__47617;
    wire N__47616;
    wire N__47615;
    wire N__47614;
    wire N__47613;
    wire N__47612;
    wire N__47611;
    wire N__47610;
    wire N__47609;
    wire N__47608;
    wire N__47607;
    wire N__47606;
    wire N__47605;
    wire N__47604;
    wire N__47603;
    wire N__47602;
    wire N__47601;
    wire N__47600;
    wire N__47599;
    wire N__47598;
    wire N__47597;
    wire N__47596;
    wire N__47595;
    wire N__47594;
    wire N__47593;
    wire N__47592;
    wire N__47591;
    wire N__47590;
    wire N__47589;
    wire N__47588;
    wire N__47587;
    wire N__47586;
    wire N__47585;
    wire N__47584;
    wire N__47583;
    wire N__47582;
    wire N__47581;
    wire N__47580;
    wire N__47579;
    wire N__47578;
    wire N__47577;
    wire N__47576;
    wire N__47575;
    wire N__47574;
    wire N__47573;
    wire N__47572;
    wire N__47571;
    wire N__47570;
    wire N__47569;
    wire N__47568;
    wire N__47567;
    wire N__47566;
    wire N__47565;
    wire N__47564;
    wire N__47563;
    wire N__47562;
    wire N__47561;
    wire N__47560;
    wire N__47559;
    wire N__47558;
    wire N__47557;
    wire N__47556;
    wire N__47555;
    wire N__47554;
    wire N__47553;
    wire N__47552;
    wire N__47551;
    wire N__47550;
    wire N__47549;
    wire N__47240;
    wire N__47237;
    wire N__47236;
    wire N__47233;
    wire N__47230;
    wire N__47229;
    wire N__47224;
    wire N__47221;
    wire N__47220;
    wire N__47219;
    wire N__47216;
    wire N__47213;
    wire N__47210;
    wire N__47209;
    wire N__47208;
    wire N__47205;
    wire N__47204;
    wire N__47203;
    wire N__47202;
    wire N__47195;
    wire N__47192;
    wire N__47191;
    wire N__47190;
    wire N__47189;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47179;
    wire N__47176;
    wire N__47173;
    wire N__47172;
    wire N__47171;
    wire N__47166;
    wire N__47165;
    wire N__47164;
    wire N__47163;
    wire N__47162;
    wire N__47161;
    wire N__47160;
    wire N__47159;
    wire N__47158;
    wire N__47157;
    wire N__47156;
    wire N__47155;
    wire N__47154;
    wire N__47153;
    wire N__47152;
    wire N__47151;
    wire N__47150;
    wire N__47147;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47126;
    wire N__47123;
    wire N__47120;
    wire N__47119;
    wire N__47118;
    wire N__47117;
    wire N__47116;
    wire N__47115;
    wire N__47114;
    wire N__47113;
    wire N__47110;
    wire N__47101;
    wire N__47092;
    wire N__47083;
    wire N__47074;
    wire N__47071;
    wire N__47070;
    wire N__47069;
    wire N__47068;
    wire N__47067;
    wire N__47062;
    wire N__47053;
    wire N__47050;
    wire N__47043;
    wire N__47034;
    wire N__47029;
    wire N__47026;
    wire N__47019;
    wire N__47010;
    wire N__47005;
    wire N__46998;
    wire N__46993;
    wire N__46990;
    wire N__46987;
    wire N__46984;
    wire N__46981;
    wire N__46978;
    wire N__46975;
    wire N__46970;
    wire N__46961;
    wire N__46960;
    wire N__46959;
    wire N__46958;
    wire N__46955;
    wire N__46950;
    wire N__46947;
    wire N__46944;
    wire N__46941;
    wire N__46940;
    wire N__46939;
    wire N__46938;
    wire N__46937;
    wire N__46936;
    wire N__46933;
    wire N__46932;
    wire N__46931;
    wire N__46930;
    wire N__46929;
    wire N__46928;
    wire N__46927;
    wire N__46926;
    wire N__46925;
    wire N__46924;
    wire N__46923;
    wire N__46922;
    wire N__46921;
    wire N__46920;
    wire N__46919;
    wire N__46918;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46913;
    wire N__46912;
    wire N__46911;
    wire N__46910;
    wire N__46909;
    wire N__46908;
    wire N__46907;
    wire N__46906;
    wire N__46905;
    wire N__46904;
    wire N__46903;
    wire N__46902;
    wire N__46901;
    wire N__46900;
    wire N__46899;
    wire N__46898;
    wire N__46897;
    wire N__46896;
    wire N__46895;
    wire N__46894;
    wire N__46893;
    wire N__46892;
    wire N__46891;
    wire N__46890;
    wire N__46889;
    wire N__46888;
    wire N__46887;
    wire N__46886;
    wire N__46885;
    wire N__46884;
    wire N__46883;
    wire N__46882;
    wire N__46881;
    wire N__46880;
    wire N__46879;
    wire N__46878;
    wire N__46877;
    wire N__46876;
    wire N__46875;
    wire N__46874;
    wire N__46873;
    wire N__46872;
    wire N__46871;
    wire N__46870;
    wire N__46869;
    wire N__46868;
    wire N__46867;
    wire N__46866;
    wire N__46865;
    wire N__46864;
    wire N__46863;
    wire N__46862;
    wire N__46861;
    wire N__46860;
    wire N__46859;
    wire N__46858;
    wire N__46857;
    wire N__46856;
    wire N__46855;
    wire N__46854;
    wire N__46853;
    wire N__46852;
    wire N__46851;
    wire N__46850;
    wire N__46849;
    wire N__46848;
    wire N__46847;
    wire N__46846;
    wire N__46845;
    wire N__46844;
    wire N__46843;
    wire N__46842;
    wire N__46841;
    wire N__46840;
    wire N__46839;
    wire N__46838;
    wire N__46837;
    wire N__46836;
    wire N__46835;
    wire N__46834;
    wire N__46833;
    wire N__46832;
    wire N__46831;
    wire N__46830;
    wire N__46829;
    wire N__46828;
    wire N__46827;
    wire N__46826;
    wire N__46825;
    wire N__46824;
    wire N__46823;
    wire N__46822;
    wire N__46821;
    wire N__46820;
    wire N__46819;
    wire N__46818;
    wire N__46817;
    wire N__46816;
    wire N__46815;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46811;
    wire N__46810;
    wire N__46809;
    wire N__46808;
    wire N__46807;
    wire N__46806;
    wire N__46805;
    wire N__46804;
    wire N__46803;
    wire N__46802;
    wire N__46801;
    wire N__46800;
    wire N__46799;
    wire N__46798;
    wire N__46797;
    wire N__46796;
    wire N__46795;
    wire N__46794;
    wire N__46793;
    wire N__46792;
    wire N__46791;
    wire N__46790;
    wire N__46789;
    wire N__46788;
    wire N__46787;
    wire N__46786;
    wire N__46785;
    wire N__46784;
    wire N__46783;
    wire N__46466;
    wire N__46463;
    wire N__46460;
    wire N__46457;
    wire N__46454;
    wire N__46451;
    wire N__46448;
    wire N__46445;
    wire N__46444;
    wire N__46439;
    wire N__46436;
    wire N__46435;
    wire N__46434;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46418;
    wire N__46415;
    wire N__46414;
    wire N__46411;
    wire N__46408;
    wire N__46403;
    wire N__46402;
    wire N__46399;
    wire N__46396;
    wire N__46393;
    wire N__46388;
    wire N__46387;
    wire N__46382;
    wire N__46379;
    wire N__46376;
    wire N__46373;
    wire N__46370;
    wire N__46367;
    wire N__46366;
    wire N__46365;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46351;
    wire N__46346;
    wire N__46345;
    wire N__46342;
    wire N__46339;
    wire N__46334;
    wire N__46331;
    wire N__46330;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46317;
    wire N__46314;
    wire N__46307;
    wire N__46306;
    wire N__46303;
    wire N__46300;
    wire N__46295;
    wire N__46292;
    wire N__46289;
    wire N__46286;
    wire N__46283;
    wire N__46280;
    wire N__46277;
    wire N__46274;
    wire N__46271;
    wire N__46270;
    wire N__46267;
    wire N__46264;
    wire N__46259;
    wire N__46256;
    wire N__46255;
    wire N__46254;
    wire N__46253;
    wire N__46250;
    wire N__46249;
    wire N__46248;
    wire N__46247;
    wire N__46244;
    wire N__46243;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46235;
    wire N__46234;
    wire N__46233;
    wire N__46232;
    wire N__46231;
    wire N__46228;
    wire N__46219;
    wire N__46210;
    wire N__46209;
    wire N__46208;
    wire N__46203;
    wire N__46196;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46184;
    wire N__46183;
    wire N__46182;
    wire N__46181;
    wire N__46180;
    wire N__46179;
    wire N__46178;
    wire N__46177;
    wire N__46176;
    wire N__46175;
    wire N__46174;
    wire N__46173;
    wire N__46172;
    wire N__46171;
    wire N__46170;
    wire N__46169;
    wire N__46166;
    wire N__46163;
    wire N__46160;
    wire N__46155;
    wire N__46152;
    wire N__46135;
    wire N__46120;
    wire N__46117;
    wire N__46114;
    wire N__46111;
    wire N__46108;
    wire N__46105;
    wire N__46098;
    wire N__46089;
    wire N__46082;
    wire N__46079;
    wire N__46076;
    wire N__46075;
    wire N__46074;
    wire N__46073;
    wire N__46072;
    wire N__46071;
    wire N__46068;
    wire N__46065;
    wire N__46064;
    wire N__46061;
    wire N__46058;
    wire N__46057;
    wire N__46054;
    wire N__46051;
    wire N__46048;
    wire N__46045;
    wire N__46038;
    wire N__46031;
    wire N__46028;
    wire N__46021;
    wire N__46018;
    wire N__46015;
    wire N__46010;
    wire N__46007;
    wire N__46004;
    wire N__46001;
    wire N__45998;
    wire N__45995;
    wire N__45992;
    wire N__45991;
    wire N__45986;
    wire N__45983;
    wire N__45980;
    wire N__45979;
    wire N__45974;
    wire N__45971;
    wire N__45970;
    wire N__45967;
    wire N__45964;
    wire N__45959;
    wire N__45958;
    wire N__45957;
    wire N__45956;
    wire N__45955;
    wire N__45954;
    wire N__45953;
    wire N__45952;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45928;
    wire N__45927;
    wire N__45926;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45914;
    wire N__45911;
    wire N__45906;
    wire N__45903;
    wire N__45900;
    wire N__45895;
    wire N__45892;
    wire N__45889;
    wire N__45884;
    wire N__45883;
    wire N__45882;
    wire N__45879;
    wire N__45876;
    wire N__45873;
    wire N__45868;
    wire N__45863;
    wire N__45862;
    wire N__45859;
    wire N__45858;
    wire N__45855;
    wire N__45852;
    wire N__45849;
    wire N__45842;
    wire N__45841;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45815;
    wire N__45812;
    wire N__45809;
    wire N__45806;
    wire N__45803;
    wire N__45800;
    wire N__45797;
    wire N__45788;
    wire N__45787;
    wire N__45786;
    wire N__45783;
    wire N__45780;
    wire N__45777;
    wire N__45770;
    wire N__45769;
    wire N__45766;
    wire N__45763;
    wire N__45758;
    wire N__45757;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45742;
    wire N__45739;
    wire N__45736;
    wire N__45731;
    wire N__45728;
    wire N__45725;
    wire N__45722;
    wire N__45719;
    wire N__45716;
    wire N__45713;
    wire N__45712;
    wire N__45709;
    wire N__45706;
    wire N__45705;
    wire N__45704;
    wire N__45699;
    wire N__45696;
    wire N__45693;
    wire N__45688;
    wire N__45685;
    wire N__45682;
    wire N__45679;
    wire N__45676;
    wire N__45673;
    wire N__45668;
    wire N__45667;
    wire N__45664;
    wire N__45663;
    wire N__45660;
    wire N__45657;
    wire N__45654;
    wire N__45647;
    wire N__45644;
    wire N__45641;
    wire N__45638;
    wire N__45637;
    wire N__45632;
    wire N__45629;
    wire N__45628;
    wire N__45623;
    wire N__45620;
    wire N__45619;
    wire N__45616;
    wire N__45615;
    wire N__45610;
    wire N__45607;
    wire N__45604;
    wire N__45599;
    wire N__45598;
    wire N__45595;
    wire N__45594;
    wire N__45589;
    wire N__45586;
    wire N__45583;
    wire N__45578;
    wire N__45575;
    wire N__45572;
    wire N__45569;
    wire N__45566;
    wire N__45563;
    wire N__45560;
    wire N__45557;
    wire N__45556;
    wire N__45555;
    wire N__45552;
    wire N__45549;
    wire N__45546;
    wire N__45543;
    wire N__45540;
    wire N__45539;
    wire N__45536;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45513;
    wire N__45506;
    wire N__45503;
    wire N__45500;
    wire N__45499;
    wire N__45498;
    wire N__45497;
    wire N__45494;
    wire N__45489;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45479;
    wire N__45476;
    wire N__45473;
    wire N__45470;
    wire N__45467;
    wire N__45462;
    wire N__45457;
    wire N__45454;
    wire N__45449;
    wire N__45448;
    wire N__45445;
    wire N__45440;
    wire N__45437;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45422;
    wire N__45419;
    wire N__45418;
    wire N__45415;
    wire N__45412;
    wire N__45407;
    wire N__45406;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45392;
    wire N__45389;
    wire N__45386;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45374;
    wire N__45371;
    wire N__45370;
    wire N__45365;
    wire N__45362;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45347;
    wire N__45346;
    wire N__45343;
    wire N__45338;
    wire N__45337;
    wire N__45334;
    wire N__45331;
    wire N__45328;
    wire N__45323;
    wire N__45320;
    wire N__45317;
    wire N__45314;
    wire N__45311;
    wire N__45310;
    wire N__45305;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45293;
    wire N__45290;
    wire N__45287;
    wire N__45286;
    wire N__45281;
    wire N__45278;
    wire N__45277;
    wire N__45276;
    wire N__45273;
    wire N__45270;
    wire N__45267;
    wire N__45262;
    wire N__45257;
    wire N__45256;
    wire N__45253;
    wire N__45250;
    wire N__45247;
    wire N__45244;
    wire N__45243;
    wire N__45238;
    wire N__45235;
    wire N__45232;
    wire N__45227;
    wire N__45226;
    wire N__45221;
    wire N__45218;
    wire N__45217;
    wire N__45212;
    wire N__45211;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45199;
    wire N__45194;
    wire N__45191;
    wire N__45190;
    wire N__45187;
    wire N__45186;
    wire N__45183;
    wire N__45182;
    wire N__45179;
    wire N__45172;
    wire N__45167;
    wire N__45166;
    wire N__45163;
    wire N__45158;
    wire N__45157;
    wire N__45154;
    wire N__45151;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45141;
    wire N__45136;
    wire N__45131;
    wire N__45128;
    wire N__45125;
    wire N__45122;
    wire N__45119;
    wire N__45116;
    wire N__45113;
    wire N__45110;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45100;
    wire N__45095;
    wire N__45092;
    wire N__45089;
    wire N__45088;
    wire N__45083;
    wire N__45080;
    wire N__45079;
    wire N__45076;
    wire N__45073;
    wire N__45072;
    wire N__45071;
    wire N__45066;
    wire N__45061;
    wire N__45056;
    wire N__45055;
    wire N__45054;
    wire N__45053;
    wire N__45052;
    wire N__45051;
    wire N__45050;
    wire N__45047;
    wire N__45046;
    wire N__45045;
    wire N__45044;
    wire N__45043;
    wire N__45040;
    wire N__45039;
    wire N__45038;
    wire N__45037;
    wire N__45036;
    wire N__45035;
    wire N__45034;
    wire N__45033;
    wire N__45032;
    wire N__45031;
    wire N__45030;
    wire N__45029;
    wire N__45028;
    wire N__45027;
    wire N__45024;
    wire N__45023;
    wire N__45020;
    wire N__45019;
    wire N__45016;
    wire N__45015;
    wire N__45014;
    wire N__45013;
    wire N__45012;
    wire N__45011;
    wire N__45010;
    wire N__45009;
    wire N__45008;
    wire N__45007;
    wire N__45006;
    wire N__45005;
    wire N__45004;
    wire N__45003;
    wire N__45000;
    wire N__44999;
    wire N__44998;
    wire N__44997;
    wire N__44996;
    wire N__44995;
    wire N__44994;
    wire N__44989;
    wire N__44986;
    wire N__44983;
    wire N__44980;
    wire N__44979;
    wire N__44976;
    wire N__44975;
    wire N__44974;
    wire N__44973;
    wire N__44972;
    wire N__44971;
    wire N__44970;
    wire N__44969;
    wire N__44966;
    wire N__44965;
    wire N__44962;
    wire N__44961;
    wire N__44958;
    wire N__44955;
    wire N__44954;
    wire N__44949;
    wire N__44948;
    wire N__44939;
    wire N__44938;
    wire N__44937;
    wire N__44936;
    wire N__44935;
    wire N__44934;
    wire N__44933;
    wire N__44932;
    wire N__44931;
    wire N__44928;
    wire N__44927;
    wire N__44926;
    wire N__44925;
    wire N__44924;
    wire N__44923;
    wire N__44920;
    wire N__44919;
    wire N__44902;
    wire N__44899;
    wire N__44898;
    wire N__44895;
    wire N__44894;
    wire N__44891;
    wire N__44890;
    wire N__44887;
    wire N__44886;
    wire N__44883;
    wire N__44882;
    wire N__44879;
    wire N__44878;
    wire N__44875;
    wire N__44874;
    wire N__44871;
    wire N__44870;
    wire N__44867;
    wire N__44866;
    wire N__44863;
    wire N__44862;
    wire N__44859;
    wire N__44858;
    wire N__44853;
    wire N__44852;
    wire N__44851;
    wire N__44850;
    wire N__44847;
    wire N__44844;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44834;
    wire N__44833;
    wire N__44830;
    wire N__44829;
    wire N__44828;
    wire N__44827;
    wire N__44824;
    wire N__44821;
    wire N__44818;
    wire N__44811;
    wire N__44810;
    wire N__44807;
    wire N__44806;
    wire N__44803;
    wire N__44802;
    wire N__44799;
    wire N__44798;
    wire N__44795;
    wire N__44794;
    wire N__44791;
    wire N__44790;
    wire N__44787;
    wire N__44786;
    wire N__44783;
    wire N__44782;
    wire N__44781;
    wire N__44780;
    wire N__44779;
    wire N__44778;
    wire N__44777;
    wire N__44776;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44764;
    wire N__44761;
    wire N__44756;
    wire N__44753;
    wire N__44750;
    wire N__44747;
    wire N__44732;
    wire N__44717;
    wire N__44712;
    wire N__44709;
    wire N__44692;
    wire N__44675;
    wire N__44662;
    wire N__44659;
    wire N__44652;
    wire N__44645;
    wire N__44628;
    wire N__44627;
    wire N__44626;
    wire N__44625;
    wire N__44624;
    wire N__44623;
    wire N__44622;
    wire N__44619;
    wire N__44612;
    wire N__44597;
    wire N__44580;
    wire N__44577;
    wire N__44576;
    wire N__44573;
    wire N__44572;
    wire N__44569;
    wire N__44568;
    wire N__44565;
    wire N__44564;
    wire N__44561;
    wire N__44560;
    wire N__44557;
    wire N__44556;
    wire N__44553;
    wire N__44552;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44518;
    wire N__44515;
    wire N__44508;
    wire N__44505;
    wire N__44494;
    wire N__44485;
    wire N__44468;
    wire N__44455;
    wire N__44446;
    wire N__44429;
    wire N__44428;
    wire N__44427;
    wire N__44426;
    wire N__44425;
    wire N__44424;
    wire N__44423;
    wire N__44422;
    wire N__44421;
    wire N__44420;
    wire N__44419;
    wire N__44418;
    wire N__44417;
    wire N__44416;
    wire N__44415;
    wire N__44414;
    wire N__44411;
    wire N__44408;
    wire N__44407;
    wire N__44406;
    wire N__44405;
    wire N__44404;
    wire N__44403;
    wire N__44402;
    wire N__44401;
    wire N__44400;
    wire N__44399;
    wire N__44398;
    wire N__44397;
    wire N__44396;
    wire N__44395;
    wire N__44394;
    wire N__44393;
    wire N__44392;
    wire N__44391;
    wire N__44390;
    wire N__44389;
    wire N__44388;
    wire N__44385;
    wire N__44382;
    wire N__44369;
    wire N__44366;
    wire N__44365;
    wire N__44364;
    wire N__44363;
    wire N__44362;
    wire N__44361;
    wire N__44360;
    wire N__44359;
    wire N__44356;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44344;
    wire N__44339;
    wire N__44336;
    wire N__44323;
    wire N__44316;
    wire N__44311;
    wire N__44302;
    wire N__44299;
    wire N__44298;
    wire N__44297;
    wire N__44296;
    wire N__44295;
    wire N__44294;
    wire N__44293;
    wire N__44292;
    wire N__44291;
    wire N__44288;
    wire N__44283;
    wire N__44282;
    wire N__44281;
    wire N__44280;
    wire N__44279;
    wire N__44278;
    wire N__44277;
    wire N__44272;
    wire N__44269;
    wire N__44252;
    wire N__44249;
    wire N__44246;
    wire N__44243;
    wire N__44240;
    wire N__44239;
    wire N__44236;
    wire N__44227;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44201;
    wire N__44200;
    wire N__44199;
    wire N__44198;
    wire N__44197;
    wire N__44196;
    wire N__44195;
    wire N__44194;
    wire N__44193;
    wire N__44192;
    wire N__44191;
    wire N__44190;
    wire N__44189;
    wire N__44184;
    wire N__44171;
    wire N__44162;
    wire N__44155;
    wire N__44152;
    wire N__44145;
    wire N__44138;
    wire N__44123;
    wire N__44118;
    wire N__44115;
    wire N__44110;
    wire N__44105;
    wire N__44102;
    wire N__44095;
    wire N__44078;
    wire N__44075;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44062;
    wire N__44061;
    wire N__44058;
    wire N__44055;
    wire N__44052;
    wire N__44047;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44029;
    wire N__44024;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44012;
    wire N__44009;
    wire N__44008;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43997;
    wire N__43990;
    wire N__43987;
    wire N__43982;
    wire N__43979;
    wire N__43976;
    wire N__43973;
    wire N__43970;
    wire N__43967;
    wire N__43966;
    wire N__43963;
    wire N__43960;
    wire N__43959;
    wire N__43956;
    wire N__43953;
    wire N__43950;
    wire N__43949;
    wire N__43946;
    wire N__43943;
    wire N__43940;
    wire N__43937;
    wire N__43934;
    wire N__43931;
    wire N__43928;
    wire N__43925;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43901;
    wire N__43900;
    wire N__43899;
    wire N__43896;
    wire N__43891;
    wire N__43890;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43876;
    wire N__43871;
    wire N__43868;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43855;
    wire N__43852;
    wire N__43851;
    wire N__43848;
    wire N__43847;
    wire N__43846;
    wire N__43845;
    wire N__43844;
    wire N__43843;
    wire N__43840;
    wire N__43837;
    wire N__43830;
    wire N__43827;
    wire N__43822;
    wire N__43821;
    wire N__43818;
    wire N__43811;
    wire N__43808;
    wire N__43805;
    wire N__43804;
    wire N__43799;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43760;
    wire N__43757;
    wire N__43754;
    wire N__43751;
    wire N__43750;
    wire N__43747;
    wire N__43744;
    wire N__43743;
    wire N__43740;
    wire N__43735;
    wire N__43730;
    wire N__43727;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43716;
    wire N__43711;
    wire N__43708;
    wire N__43703;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43688;
    wire N__43685;
    wire N__43684;
    wire N__43681;
    wire N__43680;
    wire N__43679;
    wire N__43676;
    wire N__43673;
    wire N__43668;
    wire N__43665;
    wire N__43660;
    wire N__43657;
    wire N__43654;
    wire N__43649;
    wire N__43646;
    wire N__43645;
    wire N__43644;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43628;
    wire N__43625;
    wire N__43622;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43594;
    wire N__43593;
    wire N__43590;
    wire N__43587;
    wire N__43584;
    wire N__43581;
    wire N__43574;
    wire N__43573;
    wire N__43572;
    wire N__43571;
    wire N__43570;
    wire N__43569;
    wire N__43568;
    wire N__43567;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43541;
    wire N__43538;
    wire N__43535;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43517;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43506;
    wire N__43501;
    wire N__43498;
    wire N__43493;
    wire N__43490;
    wire N__43487;
    wire N__43484;
    wire N__43481;
    wire N__43478;
    wire N__43475;
    wire N__43474;
    wire N__43473;
    wire N__43470;
    wire N__43467;
    wire N__43464;
    wire N__43457;
    wire N__43454;
    wire N__43451;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43424;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43412;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43396;
    wire N__43393;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43383;
    wire N__43378;
    wire N__43375;
    wire N__43370;
    wire N__43367;
    wire N__43364;
    wire N__43361;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43349;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43341;
    wire N__43338;
    wire N__43335;
    wire N__43332;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43310;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43290;
    wire N__43285;
    wire N__43282;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43232;
    wire N__43229;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43216;
    wire N__43211;
    wire N__43210;
    wire N__43207;
    wire N__43204;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43187;
    wire N__43184;
    wire N__43183;
    wire N__43178;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43148;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43140;
    wire N__43137;
    wire N__43134;
    wire N__43131;
    wire N__43124;
    wire N__43121;
    wire N__43118;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43101;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43069;
    wire N__43066;
    wire N__43063;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43046;
    wire N__43043;
    wire N__43040;
    wire N__43037;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43008;
    wire N__43001;
    wire N__42998;
    wire N__42995;
    wire N__42994;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42955;
    wire N__42952;
    wire N__42949;
    wire N__42948;
    wire N__42943;
    wire N__42940;
    wire N__42935;
    wire N__42932;
    wire N__42931;
    wire N__42928;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42910;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42896;
    wire N__42893;
    wire N__42890;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42880;
    wire N__42877;
    wire N__42876;
    wire N__42871;
    wire N__42868;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42854;
    wire N__42851;
    wire N__42848;
    wire N__42845;
    wire N__42844;
    wire N__42839;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42827;
    wire N__42824;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42799;
    wire N__42796;
    wire N__42793;
    wire N__42792;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42776;
    wire N__42773;
    wire N__42770;
    wire N__42767;
    wire N__42764;
    wire N__42761;
    wire N__42760;
    wire N__42757;
    wire N__42754;
    wire N__42751;
    wire N__42748;
    wire N__42747;
    wire N__42742;
    wire N__42739;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42725;
    wire N__42722;
    wire N__42719;
    wire N__42716;
    wire N__42715;
    wire N__42712;
    wire N__42709;
    wire N__42706;
    wire N__42703;
    wire N__42702;
    wire N__42697;
    wire N__42694;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42674;
    wire N__42671;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42660;
    wire N__42655;
    wire N__42652;
    wire N__42647;
    wire N__42644;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42631;
    wire N__42628;
    wire N__42625;
    wire N__42622;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42605;
    wire N__42602;
    wire N__42599;
    wire N__42598;
    wire N__42597;
    wire N__42596;
    wire N__42593;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42560;
    wire N__42559;
    wire N__42554;
    wire N__42551;
    wire N__42548;
    wire N__42547;
    wire N__42546;
    wire N__42545;
    wire N__42542;
    wire N__42537;
    wire N__42534;
    wire N__42529;
    wire N__42526;
    wire N__42523;
    wire N__42518;
    wire N__42517;
    wire N__42514;
    wire N__42511;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42488;
    wire N__42485;
    wire N__42482;
    wire N__42479;
    wire N__42476;
    wire N__42473;
    wire N__42470;
    wire N__42467;
    wire N__42466;
    wire N__42463;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42445;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42435;
    wire N__42428;
    wire N__42425;
    wire N__42422;
    wire N__42419;
    wire N__42416;
    wire N__42415;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42400;
    wire N__42397;
    wire N__42394;
    wire N__42391;
    wire N__42388;
    wire N__42383;
    wire N__42382;
    wire N__42381;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42370;
    wire N__42369;
    wire N__42368;
    wire N__42367;
    wire N__42366;
    wire N__42365;
    wire N__42364;
    wire N__42363;
    wire N__42362;
    wire N__42361;
    wire N__42360;
    wire N__42359;
    wire N__42358;
    wire N__42355;
    wire N__42352;
    wire N__42349;
    wire N__42346;
    wire N__42331;
    wire N__42318;
    wire N__42317;
    wire N__42316;
    wire N__42315;
    wire N__42314;
    wire N__42313;
    wire N__42312;
    wire N__42311;
    wire N__42310;
    wire N__42305;
    wire N__42296;
    wire N__42287;
    wire N__42278;
    wire N__42275;
    wire N__42266;
    wire N__42265;
    wire N__42262;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42247;
    wire N__42242;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42227;
    wire N__42226;
    wire N__42221;
    wire N__42218;
    wire N__42217;
    wire N__42214;
    wire N__42211;
    wire N__42206;
    wire N__42203;
    wire N__42200;
    wire N__42197;
    wire N__42194;
    wire N__42191;
    wire N__42190;
    wire N__42187;
    wire N__42184;
    wire N__42181;
    wire N__42178;
    wire N__42177;
    wire N__42172;
    wire N__42169;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42152;
    wire N__42149;
    wire N__42146;
    wire N__42145;
    wire N__42142;
    wire N__42139;
    wire N__42136;
    wire N__42133;
    wire N__42130;
    wire N__42127;
    wire N__42122;
    wire N__42121;
    wire N__42118;
    wire N__42115;
    wire N__42110;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42100;
    wire N__42097;
    wire N__42094;
    wire N__42091;
    wire N__42086;
    wire N__42083;
    wire N__42080;
    wire N__42077;
    wire N__42074;
    wire N__42071;
    wire N__42068;
    wire N__42065;
    wire N__42062;
    wire N__42059;
    wire N__42058;
    wire N__42055;
    wire N__42052;
    wire N__42047;
    wire N__42044;
    wire N__42041;
    wire N__42040;
    wire N__42037;
    wire N__42034;
    wire N__42031;
    wire N__42028;
    wire N__42025;
    wire N__42022;
    wire N__42021;
    wire N__42020;
    wire N__42017;
    wire N__42014;
    wire N__42009;
    wire N__42002;
    wire N__41999;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41987;
    wire N__41984;
    wire N__41983;
    wire N__41982;
    wire N__41979;
    wire N__41974;
    wire N__41969;
    wire N__41968;
    wire N__41965;
    wire N__41964;
    wire N__41961;
    wire N__41956;
    wire N__41951;
    wire N__41948;
    wire N__41945;
    wire N__41942;
    wire N__41939;
    wire N__41936;
    wire N__41935;
    wire N__41932;
    wire N__41929;
    wire N__41926;
    wire N__41925;
    wire N__41922;
    wire N__41919;
    wire N__41916;
    wire N__41911;
    wire N__41906;
    wire N__41905;
    wire N__41904;
    wire N__41901;
    wire N__41900;
    wire N__41897;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41885;
    wire N__41880;
    wire N__41877;
    wire N__41872;
    wire N__41867;
    wire N__41864;
    wire N__41863;
    wire N__41858;
    wire N__41855;
    wire N__41852;
    wire N__41849;
    wire N__41846;
    wire N__41845;
    wire N__41842;
    wire N__41839;
    wire N__41834;
    wire N__41833;
    wire N__41830;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41813;
    wire N__41810;
    wire N__41809;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41792;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41780;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41765;
    wire N__41764;
    wire N__41761;
    wire N__41758;
    wire N__41755;
    wire N__41754;
    wire N__41749;
    wire N__41746;
    wire N__41741;
    wire N__41740;
    wire N__41739;
    wire N__41738;
    wire N__41735;
    wire N__41732;
    wire N__41729;
    wire N__41726;
    wire N__41723;
    wire N__41720;
    wire N__41717;
    wire N__41712;
    wire N__41707;
    wire N__41704;
    wire N__41701;
    wire N__41698;
    wire N__41693;
    wire N__41692;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41675;
    wire N__41674;
    wire N__41673;
    wire N__41672;
    wire N__41669;
    wire N__41666;
    wire N__41663;
    wire N__41660;
    wire N__41657;
    wire N__41652;
    wire N__41649;
    wire N__41644;
    wire N__41641;
    wire N__41638;
    wire N__41635;
    wire N__41630;
    wire N__41629;
    wire N__41626;
    wire N__41623;
    wire N__41618;
    wire N__41615;
    wire N__41612;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41602;
    wire N__41597;
    wire N__41594;
    wire N__41593;
    wire N__41588;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41573;
    wire N__41572;
    wire N__41569;
    wire N__41568;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41552;
    wire N__41551;
    wire N__41548;
    wire N__41543;
    wire N__41540;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41528;
    wire N__41525;
    wire N__41524;
    wire N__41521;
    wire N__41520;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41504;
    wire N__41503;
    wire N__41502;
    wire N__41501;
    wire N__41498;
    wire N__41495;
    wire N__41492;
    wire N__41489;
    wire N__41484;
    wire N__41479;
    wire N__41474;
    wire N__41471;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41459;
    wire N__41456;
    wire N__41455;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41447;
    wire N__41444;
    wire N__41439;
    wire N__41436;
    wire N__41433;
    wire N__41428;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41416;
    wire N__41415;
    wire N__41412;
    wire N__41409;
    wire N__41406;
    wire N__41401;
    wire N__41396;
    wire N__41395;
    wire N__41394;
    wire N__41389;
    wire N__41386;
    wire N__41383;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41371;
    wire N__41368;
    wire N__41365;
    wire N__41362;
    wire N__41357;
    wire N__41354;
    wire N__41353;
    wire N__41352;
    wire N__41351;
    wire N__41350;
    wire N__41349;
    wire N__41348;
    wire N__41347;
    wire N__41346;
    wire N__41345;
    wire N__41344;
    wire N__41343;
    wire N__41342;
    wire N__41341;
    wire N__41340;
    wire N__41339;
    wire N__41338;
    wire N__41337;
    wire N__41336;
    wire N__41335;
    wire N__41334;
    wire N__41333;
    wire N__41332;
    wire N__41331;
    wire N__41330;
    wire N__41329;
    wire N__41328;
    wire N__41327;
    wire N__41326;
    wire N__41325;
    wire N__41316;
    wire N__41307;
    wire N__41302;
    wire N__41293;
    wire N__41284;
    wire N__41275;
    wire N__41266;
    wire N__41257;
    wire N__41254;
    wire N__41247;
    wire N__41240;
    wire N__41237;
    wire N__41234;
    wire N__41229;
    wire N__41224;
    wire N__41219;
    wire N__41216;
    wire N__41213;
    wire N__41212;
    wire N__41209;
    wire N__41206;
    wire N__41203;
    wire N__41198;
    wire N__41197;
    wire N__41194;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41163;
    wire N__41160;
    wire N__41155;
    wire N__41150;
    wire N__41149;
    wire N__41148;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41136;
    wire N__41133;
    wire N__41128;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41114;
    wire N__41113;
    wire N__41112;
    wire N__41111;
    wire N__41106;
    wire N__41103;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41091;
    wire N__41088;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41076;
    wire N__41069;
    wire N__41066;
    wire N__41063;
    wire N__41062;
    wire N__41059;
    wire N__41056;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41046;
    wire N__41045;
    wire N__41042;
    wire N__41039;
    wire N__41034;
    wire N__41031;
    wire N__41024;
    wire N__41021;
    wire N__41018;
    wire N__41017;
    wire N__41016;
    wire N__41011;
    wire N__41008;
    wire N__41005;
    wire N__41000;
    wire N__40997;
    wire N__40994;
    wire N__40993;
    wire N__40992;
    wire N__40989;
    wire N__40986;
    wire N__40983;
    wire N__40978;
    wire N__40973;
    wire N__40970;
    wire N__40969;
    wire N__40966;
    wire N__40963;
    wire N__40962;
    wire N__40957;
    wire N__40954;
    wire N__40951;
    wire N__40946;
    wire N__40943;
    wire N__40942;
    wire N__40941;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40925;
    wire N__40922;
    wire N__40921;
    wire N__40920;
    wire N__40915;
    wire N__40912;
    wire N__40909;
    wire N__40904;
    wire N__40901;
    wire N__40900;
    wire N__40897;
    wire N__40894;
    wire N__40893;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40877;
    wire N__40874;
    wire N__40873;
    wire N__40870;
    wire N__40867;
    wire N__40864;
    wire N__40863;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40841;
    wire N__40838;
    wire N__40837;
    wire N__40834;
    wire N__40831;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40815;
    wire N__40808;
    wire N__40805;
    wire N__40804;
    wire N__40803;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40787;
    wire N__40784;
    wire N__40783;
    wire N__40782;
    wire N__40777;
    wire N__40774;
    wire N__40771;
    wire N__40766;
    wire N__40763;
    wire N__40762;
    wire N__40761;
    wire N__40756;
    wire N__40753;
    wire N__40750;
    wire N__40745;
    wire N__40742;
    wire N__40741;
    wire N__40738;
    wire N__40737;
    wire N__40734;
    wire N__40731;
    wire N__40728;
    wire N__40723;
    wire N__40718;
    wire N__40715;
    wire N__40714;
    wire N__40711;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40701;
    wire N__40696;
    wire N__40691;
    wire N__40688;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40680;
    wire N__40675;
    wire N__40672;
    wire N__40669;
    wire N__40664;
    wire N__40661;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40653;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40637;
    wire N__40634;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40604;
    wire N__40601;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40587;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40571;
    wire N__40568;
    wire N__40567;
    wire N__40566;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40550;
    wire N__40547;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40536;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40520;
    wire N__40517;
    wire N__40516;
    wire N__40513;
    wire N__40510;
    wire N__40509;
    wire N__40504;
    wire N__40501;
    wire N__40498;
    wire N__40493;
    wire N__40490;
    wire N__40489;
    wire N__40486;
    wire N__40483;
    wire N__40482;
    wire N__40477;
    wire N__40474;
    wire N__40471;
    wire N__40466;
    wire N__40463;
    wire N__40462;
    wire N__40461;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40445;
    wire N__40442;
    wire N__40441;
    wire N__40440;
    wire N__40435;
    wire N__40432;
    wire N__40429;
    wire N__40424;
    wire N__40421;
    wire N__40420;
    wire N__40417;
    wire N__40414;
    wire N__40413;
    wire N__40410;
    wire N__40407;
    wire N__40404;
    wire N__40399;
    wire N__40394;
    wire N__40391;
    wire N__40388;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40360;
    wire N__40355;
    wire N__40352;
    wire N__40349;
    wire N__40348;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40328;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40310;
    wire N__40307;
    wire N__40304;
    wire N__40303;
    wire N__40302;
    wire N__40297;
    wire N__40294;
    wire N__40289;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40277;
    wire N__40274;
    wire N__40271;
    wire N__40268;
    wire N__40265;
    wire N__40262;
    wire N__40261;
    wire N__40260;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40239;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40220;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40202;
    wire N__40199;
    wire N__40196;
    wire N__40193;
    wire N__40192;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40178;
    wire N__40175;
    wire N__40170;
    wire N__40167;
    wire N__40160;
    wire N__40157;
    wire N__40154;
    wire N__40153;
    wire N__40150;
    wire N__40147;
    wire N__40146;
    wire N__40143;
    wire N__40140;
    wire N__40137;
    wire N__40132;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40120;
    wire N__40117;
    wire N__40114;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40096;
    wire N__40095;
    wire N__40090;
    wire N__40087;
    wire N__40082;
    wire N__40079;
    wire N__40076;
    wire N__40073;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40065;
    wire N__40062;
    wire N__40059;
    wire N__40056;
    wire N__40053;
    wire N__40052;
    wire N__40049;
    wire N__40046;
    wire N__40043;
    wire N__40040;
    wire N__40031;
    wire N__40028;
    wire N__40025;
    wire N__40022;
    wire N__40019;
    wire N__40018;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40003;
    wire N__40000;
    wire N__39999;
    wire N__39994;
    wire N__39991;
    wire N__39986;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39974;
    wire N__39971;
    wire N__39970;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39952;
    wire N__39951;
    wire N__39946;
    wire N__39943;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39929;
    wire N__39926;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39904;
    wire N__39901;
    wire N__39900;
    wire N__39895;
    wire N__39892;
    wire N__39887;
    wire N__39884;
    wire N__39881;
    wire N__39878;
    wire N__39877;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39860;
    wire N__39857;
    wire N__39852;
    wire N__39849;
    wire N__39842;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39823;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39813;
    wire N__39808;
    wire N__39805;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39795;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39764;
    wire N__39761;
    wire N__39758;
    wire N__39757;
    wire N__39754;
    wire N__39751;
    wire N__39750;
    wire N__39747;
    wire N__39744;
    wire N__39741;
    wire N__39736;
    wire N__39733;
    wire N__39728;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39716;
    wire N__39713;
    wire N__39710;
    wire N__39709;
    wire N__39706;
    wire N__39703;
    wire N__39702;
    wire N__39697;
    wire N__39694;
    wire N__39691;
    wire N__39688;
    wire N__39687;
    wire N__39682;
    wire N__39679;
    wire N__39674;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39664;
    wire N__39661;
    wire N__39660;
    wire N__39657;
    wire N__39654;
    wire N__39651;
    wire N__39648;
    wire N__39643;
    wire N__39642;
    wire N__39637;
    wire N__39634;
    wire N__39629;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39619;
    wire N__39616;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39603;
    wire N__39600;
    wire N__39597;
    wire N__39596;
    wire N__39593;
    wire N__39588;
    wire N__39585;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39571;
    wire N__39568;
    wire N__39567;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39553;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39536;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39526;
    wire N__39525;
    wire N__39522;
    wire N__39517;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39494;
    wire N__39493;
    wire N__39490;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39475;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39448;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39434;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39416;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39406;
    wire N__39405;
    wire N__39400;
    wire N__39397;
    wire N__39392;
    wire N__39391;
    wire N__39388;
    wire N__39385;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39373;
    wire N__39370;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39351;
    wire N__39350;
    wire N__39343;
    wire N__39340;
    wire N__39335;
    wire N__39332;
    wire N__39329;
    wire N__39326;
    wire N__39325;
    wire N__39322;
    wire N__39321;
    wire N__39316;
    wire N__39313;
    wire N__39310;
    wire N__39307;
    wire N__39306;
    wire N__39301;
    wire N__39298;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39284;
    wire N__39281;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39266;
    wire N__39263;
    wire N__39258;
    wire N__39255;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39239;
    wire N__39236;
    wire N__39235;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39220;
    wire N__39215;
    wire N__39212;
    wire N__39209;
    wire N__39208;
    wire N__39207;
    wire N__39202;
    wire N__39199;
    wire N__39196;
    wire N__39191;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39179;
    wire N__39176;
    wire N__39173;
    wire N__39170;
    wire N__39169;
    wire N__39166;
    wire N__39165;
    wire N__39160;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39137;
    wire N__39134;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39122;
    wire N__39119;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39107;
    wire N__39104;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39092;
    wire N__39089;
    wire N__39086;
    wire N__39083;
    wire N__39080;
    wire N__39077;
    wire N__39076;
    wire N__39073;
    wire N__39072;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39056;
    wire N__39053;
    wire N__39052;
    wire N__39051;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39035;
    wire N__39032;
    wire N__39031;
    wire N__39028;
    wire N__39025;
    wire N__39020;
    wire N__39017;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39005;
    wire N__39002;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38990;
    wire N__38987;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38975;
    wire N__38972;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38960;
    wire N__38957;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38945;
    wire N__38942;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38930;
    wire N__38927;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38915;
    wire N__38912;
    wire N__38911;
    wire N__38910;
    wire N__38907;
    wire N__38904;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38888;
    wire N__38885;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38867;
    wire N__38866;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38851;
    wire N__38846;
    wire N__38843;
    wire N__38842;
    wire N__38841;
    wire N__38838;
    wire N__38833;
    wire N__38830;
    wire N__38825;
    wire N__38824;
    wire N__38821;
    wire N__38818;
    wire N__38817;
    wire N__38814;
    wire N__38809;
    wire N__38806;
    wire N__38801;
    wire N__38798;
    wire N__38797;
    wire N__38796;
    wire N__38795;
    wire N__38792;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38773;
    wire N__38770;
    wire N__38767;
    wire N__38762;
    wire N__38759;
    wire N__38758;
    wire N__38755;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38738;
    wire N__38737;
    wire N__38736;
    wire N__38735;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38699;
    wire N__38698;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38674;
    wire N__38671;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38653;
    wire N__38648;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38636;
    wire N__38633;
    wire N__38632;
    wire N__38629;
    wire N__38626;
    wire N__38621;
    wire N__38618;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38594;
    wire N__38591;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38579;
    wire N__38576;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38564;
    wire N__38561;
    wire N__38558;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38546;
    wire N__38543;
    wire N__38542;
    wire N__38537;
    wire N__38534;
    wire N__38531;
    wire N__38528;
    wire N__38525;
    wire N__38522;
    wire N__38521;
    wire N__38520;
    wire N__38517;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38501;
    wire N__38500;
    wire N__38499;
    wire N__38498;
    wire N__38495;
    wire N__38490;
    wire N__38487;
    wire N__38482;
    wire N__38479;
    wire N__38476;
    wire N__38471;
    wire N__38468;
    wire N__38465;
    wire N__38462;
    wire N__38459;
    wire N__38458;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38444;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38428;
    wire N__38423;
    wire N__38420;
    wire N__38417;
    wire N__38414;
    wire N__38413;
    wire N__38410;
    wire N__38407;
    wire N__38402;
    wire N__38399;
    wire N__38396;
    wire N__38395;
    wire N__38390;
    wire N__38387;
    wire N__38384;
    wire N__38381;
    wire N__38378;
    wire N__38375;
    wire N__38372;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38344;
    wire N__38343;
    wire N__38342;
    wire N__38339;
    wire N__38336;
    wire N__38331;
    wire N__38328;
    wire N__38321;
    wire N__38318;
    wire N__38315;
    wire N__38312;
    wire N__38309;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38301;
    wire N__38300;
    wire N__38295;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38272;
    wire N__38267;
    wire N__38266;
    wire N__38265;
    wire N__38264;
    wire N__38259;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38244;
    wire N__38241;
    wire N__38236;
    wire N__38231;
    wire N__38228;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38217;
    wire N__38214;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38204;
    wire N__38201;
    wire N__38192;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38170;
    wire N__38165;
    wire N__38162;
    wire N__38161;
    wire N__38160;
    wire N__38159;
    wire N__38156;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38132;
    wire N__38127;
    wire N__38120;
    wire N__38119;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38099;
    wire N__38098;
    wire N__38097;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38081;
    wire N__38080;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38060;
    wire N__38057;
    wire N__38056;
    wire N__38055;
    wire N__38050;
    wire N__38047;
    wire N__38046;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38024;
    wire N__38021;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38003;
    wire N__38002;
    wire N__38001;
    wire N__38000;
    wire N__37999;
    wire N__37998;
    wire N__37997;
    wire N__37996;
    wire N__37995;
    wire N__37994;
    wire N__37993;
    wire N__37992;
    wire N__37991;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37981;
    wire N__37980;
    wire N__37979;
    wire N__37978;
    wire N__37977;
    wire N__37976;
    wire N__37975;
    wire N__37972;
    wire N__37971;
    wire N__37968;
    wire N__37967;
    wire N__37964;
    wire N__37963;
    wire N__37960;
    wire N__37959;
    wire N__37956;
    wire N__37955;
    wire N__37952;
    wire N__37951;
    wire N__37948;
    wire N__37947;
    wire N__37944;
    wire N__37943;
    wire N__37940;
    wire N__37939;
    wire N__37936;
    wire N__37935;
    wire N__37932;
    wire N__37931;
    wire N__37930;
    wire N__37929;
    wire N__37928;
    wire N__37921;
    wire N__37918;
    wire N__37917;
    wire N__37914;
    wire N__37909;
    wire N__37906;
    wire N__37905;
    wire N__37904;
    wire N__37903;
    wire N__37902;
    wire N__37901;
    wire N__37900;
    wire N__37899;
    wire N__37898;
    wire N__37897;
    wire N__37894;
    wire N__37879;
    wire N__37864;
    wire N__37847;
    wire N__37846;
    wire N__37845;
    wire N__37844;
    wire N__37843;
    wire N__37840;
    wire N__37835;
    wire N__37830;
    wire N__37829;
    wire N__37828;
    wire N__37827;
    wire N__37826;
    wire N__37825;
    wire N__37824;
    wire N__37823;
    wire N__37822;
    wire N__37819;
    wire N__37818;
    wire N__37815;
    wire N__37810;
    wire N__37807;
    wire N__37804;
    wire N__37797;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37777;
    wire N__37774;
    wire N__37773;
    wire N__37770;
    wire N__37769;
    wire N__37766;
    wire N__37765;
    wire N__37762;
    wire N__37761;
    wire N__37760;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37743;
    wire N__37734;
    wire N__37727;
    wire N__37720;
    wire N__37711;
    wire N__37706;
    wire N__37689;
    wire N__37684;
    wire N__37679;
    wire N__37670;
    wire N__37667;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37644;
    wire N__37637;
    wire N__37634;
    wire N__37633;
    wire N__37632;
    wire N__37631;
    wire N__37628;
    wire N__37625;
    wire N__37624;
    wire N__37623;
    wire N__37622;
    wire N__37621;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37602;
    wire N__37601;
    wire N__37600;
    wire N__37599;
    wire N__37598;
    wire N__37595;
    wire N__37594;
    wire N__37593;
    wire N__37590;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37578;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37552;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37505;
    wire N__37502;
    wire N__37501;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37487;
    wire N__37484;
    wire N__37481;
    wire N__37478;
    wire N__37475;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37430;
    wire N__37427;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37394;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37358;
    wire N__37355;
    wire N__37352;
    wire N__37349;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37321;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37309;
    wire N__37306;
    wire N__37305;
    wire N__37302;
    wire N__37299;
    wire N__37296;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37282;
    wire N__37281;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37269;
    wire N__37262;
    wire N__37261;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37248;
    wire N__37247;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37235;
    wire N__37230;
    wire N__37227;
    wire N__37220;
    wire N__37217;
    wire N__37216;
    wire N__37213;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37198;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37060;
    wire N__37059;
    wire N__37058;
    wire N__37055;
    wire N__37048;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37033;
    wire N__37032;
    wire N__37031;
    wire N__37028;
    wire N__37021;
    wire N__37016;
    wire N__37015;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36976;
    wire N__36971;
    wire N__36970;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36956;
    wire N__36953;
    wire N__36952;
    wire N__36947;
    wire N__36946;
    wire N__36943;
    wire N__36940;
    wire N__36937;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36925;
    wire N__36920;
    wire N__36917;
    wire N__36914;
    wire N__36913;
    wire N__36908;
    wire N__36905;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36889;
    wire N__36888;
    wire N__36885;
    wire N__36880;
    wire N__36875;
    wire N__36872;
    wire N__36869;
    wire N__36866;
    wire N__36863;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36851;
    wire N__36848;
    wire N__36845;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36835;
    wire N__36830;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36815;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36802;
    wire N__36801;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36785;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36728;
    wire N__36725;
    wire N__36722;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36710;
    wire N__36709;
    wire N__36704;
    wire N__36703;
    wire N__36700;
    wire N__36697;
    wire N__36696;
    wire N__36695;
    wire N__36694;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36679;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36664;
    wire N__36661;
    wire N__36650;
    wire N__36649;
    wire N__36646;
    wire N__36643;
    wire N__36640;
    wire N__36637;
    wire N__36636;
    wire N__36635;
    wire N__36634;
    wire N__36631;
    wire N__36628;
    wire N__36625;
    wire N__36622;
    wire N__36619;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36587;
    wire N__36586;
    wire N__36583;
    wire N__36580;
    wire N__36579;
    wire N__36578;
    wire N__36577;
    wire N__36576;
    wire N__36571;
    wire N__36568;
    wire N__36565;
    wire N__36560;
    wire N__36555;
    wire N__36552;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36461;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36449;
    wire N__36446;
    wire N__36443;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36419;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36395;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36287;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36279;
    wire N__36276;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36257;
    wire N__36254;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36239;
    wire N__36236;
    wire N__36235;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36197;
    wire N__36194;
    wire N__36193;
    wire N__36192;
    wire N__36189;
    wire N__36186;
    wire N__36183;
    wire N__36178;
    wire N__36173;
    wire N__36170;
    wire N__36167;
    wire N__36166;
    wire N__36163;
    wire N__36160;
    wire N__36159;
    wire N__36158;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36119;
    wire N__36116;
    wire N__36113;
    wire N__36108;
    wire N__36103;
    wire N__36098;
    wire N__36095;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__36001;
    wire N__36000;
    wire N__35997;
    wire N__35994;
    wire N__35991;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35977;
    wire N__35976;
    wire N__35971;
    wire N__35968;
    wire N__35965;
    wire N__35960;
    wire N__35957;
    wire N__35956;
    wire N__35955;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35939;
    wire N__35936;
    wire N__35935;
    wire N__35932;
    wire N__35931;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35917;
    wire N__35912;
    wire N__35909;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35901;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35885;
    wire N__35882;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35874;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35851;
    wire N__35848;
    wire N__35845;
    wire N__35844;
    wire N__35839;
    wire N__35836;
    wire N__35833;
    wire N__35828;
    wire N__35825;
    wire N__35824;
    wire N__35823;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35801;
    wire N__35798;
    wire N__35795;
    wire N__35794;
    wire N__35793;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35770;
    wire N__35769;
    wire N__35766;
    wire N__35763;
    wire N__35760;
    wire N__35755;
    wire N__35750;
    wire N__35747;
    wire N__35746;
    wire N__35743;
    wire N__35740;
    wire N__35739;
    wire N__35734;
    wire N__35731;
    wire N__35728;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35716;
    wire N__35715;
    wire N__35712;
    wire N__35709;
    wire N__35706;
    wire N__35701;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35689;
    wire N__35688;
    wire N__35685;
    wire N__35682;
    wire N__35679;
    wire N__35674;
    wire N__35669;
    wire N__35666;
    wire N__35665;
    wire N__35664;
    wire N__35661;
    wire N__35656;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35644;
    wire N__35641;
    wire N__35638;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35628;
    wire N__35623;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35611;
    wire N__35608;
    wire N__35605;
    wire N__35604;
    wire N__35601;
    wire N__35598;
    wire N__35595;
    wire N__35588;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35577;
    wire N__35574;
    wire N__35571;
    wire N__35568;
    wire N__35565;
    wire N__35558;
    wire N__35555;
    wire N__35554;
    wire N__35551;
    wire N__35548;
    wire N__35547;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35531;
    wire N__35528;
    wire N__35527;
    wire N__35526;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35503;
    wire N__35502;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35488;
    wire N__35483;
    wire N__35480;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35472;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35456;
    wire N__35453;
    wire N__35452;
    wire N__35451;
    wire N__35448;
    wire N__35443;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35429;
    wire N__35428;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35413;
    wire N__35408;
    wire N__35405;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35394;
    wire N__35391;
    wire N__35388;
    wire N__35385;
    wire N__35382;
    wire N__35379;
    wire N__35372;
    wire N__35369;
    wire N__35366;
    wire N__35363;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35320;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35296;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35273;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35219;
    wire N__35216;
    wire N__35213;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35132;
    wire N__35129;
    wire N__35126;
    wire N__35123;
    wire N__35120;
    wire N__35117;
    wire N__35114;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35102;
    wire N__35099;
    wire N__35096;
    wire N__35093;
    wire N__35090;
    wire N__35087;
    wire N__35084;
    wire N__35081;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35071;
    wire N__35068;
    wire N__35065;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35033;
    wire N__35030;
    wire N__35027;
    wire N__35024;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35003;
    wire N__35000;
    wire N__34997;
    wire N__34994;
    wire N__34991;
    wire N__34988;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34976;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34936;
    wire N__34933;
    wire N__34930;
    wire N__34925;
    wire N__34922;
    wire N__34919;
    wire N__34916;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34894;
    wire N__34893;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34871;
    wire N__34868;
    wire N__34865;
    wire N__34862;
    wire N__34861;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34844;
    wire N__34843;
    wire N__34842;
    wire N__34839;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34823;
    wire N__34814;
    wire N__34811;
    wire N__34808;
    wire N__34805;
    wire N__34802;
    wire N__34801;
    wire N__34796;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34781;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34767;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34751;
    wire N__34750;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34729;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34714;
    wire N__34711;
    wire N__34708;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34694;
    wire N__34691;
    wire N__34690;
    wire N__34689;
    wire N__34688;
    wire N__34685;
    wire N__34682;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34663;
    wire N__34662;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34642;
    wire N__34637;
    wire N__34634;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34615;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34602;
    wire N__34597;
    wire N__34592;
    wire N__34589;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34574;
    wire N__34573;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34561;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34534;
    wire N__34533;
    wire N__34530;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34520;
    wire N__34517;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34496;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34481;
    wire N__34478;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34466;
    wire N__34463;
    wire N__34460;
    wire N__34457;
    wire N__34454;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34439;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34427;
    wire N__34424;
    wire N__34421;
    wire N__34418;
    wire N__34415;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34397;
    wire N__34394;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34364;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34331;
    wire N__34328;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34313;
    wire N__34310;
    wire N__34307;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34292;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34280;
    wire N__34277;
    wire N__34274;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34262;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34207;
    wire N__34206;
    wire N__34205;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34187;
    wire N__34184;
    wire N__34183;
    wire N__34182;
    wire N__34181;
    wire N__34180;
    wire N__34179;
    wire N__34178;
    wire N__34177;
    wire N__34176;
    wire N__34175;
    wire N__34174;
    wire N__34173;
    wire N__34172;
    wire N__34171;
    wire N__34170;
    wire N__34169;
    wire N__34168;
    wire N__34167;
    wire N__34166;
    wire N__34165;
    wire N__34164;
    wire N__34163;
    wire N__34162;
    wire N__34161;
    wire N__34152;
    wire N__34149;
    wire N__34148;
    wire N__34147;
    wire N__34146;
    wire N__34145;
    wire N__34144;
    wire N__34143;
    wire N__34142;
    wire N__34133;
    wire N__34126;
    wire N__34117;
    wire N__34108;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34092;
    wire N__34083;
    wire N__34076;
    wire N__34073;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34046;
    wire N__34041;
    wire N__34034;
    wire N__34031;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34023;
    wire N__34016;
    wire N__34015;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34001;
    wire N__33998;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33986;
    wire N__33983;
    wire N__33980;
    wire N__33979;
    wire N__33978;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33955;
    wire N__33954;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33889;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33847;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33791;
    wire N__33788;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33764;
    wire N__33763;
    wire N__33762;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33742;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33722;
    wire N__33719;
    wire N__33716;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33638;
    wire N__33635;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33623;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33569;
    wire N__33566;
    wire N__33563;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33545;
    wire N__33542;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33503;
    wire N__33500;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33449;
    wire N__33446;
    wire N__33445;
    wire N__33444;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33432;
    wire N__33429;
    wire N__33422;
    wire N__33421;
    wire N__33420;
    wire N__33419;
    wire N__33418;
    wire N__33417;
    wire N__33416;
    wire N__33415;
    wire N__33414;
    wire N__33413;
    wire N__33412;
    wire N__33411;
    wire N__33410;
    wire N__33409;
    wire N__33408;
    wire N__33407;
    wire N__33406;
    wire N__33405;
    wire N__33404;
    wire N__33403;
    wire N__33402;
    wire N__33401;
    wire N__33400;
    wire N__33399;
    wire N__33398;
    wire N__33397;
    wire N__33396;
    wire N__33395;
    wire N__33394;
    wire N__33393;
    wire N__33384;
    wire N__33375;
    wire N__33370;
    wire N__33361;
    wire N__33352;
    wire N__33343;
    wire N__33334;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33314;
    wire N__33305;
    wire N__33296;
    wire N__33293;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33245;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33237;
    wire N__33236;
    wire N__33233;
    wire N__33230;
    wire N__33227;
    wire N__33224;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33203;
    wire N__33200;
    wire N__33199;
    wire N__33196;
    wire N__33195;
    wire N__33194;
    wire N__33191;
    wire N__33184;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33128;
    wire N__33125;
    wire N__33122;
    wire N__33119;
    wire N__33118;
    wire N__33115;
    wire N__33114;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33079;
    wire N__33078;
    wire N__33077;
    wire N__33076;
    wire N__33073;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33057;
    wire N__33050;
    wire N__33049;
    wire N__33046;
    wire N__33043;
    wire N__33038;
    wire N__33035;
    wire N__33032;
    wire N__33029;
    wire N__33026;
    wire N__33025;
    wire N__33024;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33003;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32948;
    wire N__32947;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32927;
    wire N__32926;
    wire N__32921;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32891;
    wire N__32890;
    wire N__32887;
    wire N__32884;
    wire N__32879;
    wire N__32878;
    wire N__32875;
    wire N__32872;
    wire N__32871;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32859;
    wire N__32852;
    wire N__32851;
    wire N__32848;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32831;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32813;
    wire N__32812;
    wire N__32811;
    wire N__32808;
    wire N__32803;
    wire N__32802;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32790;
    wire N__32783;
    wire N__32780;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32741;
    wire N__32738;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32693;
    wire N__32690;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32671;
    wire N__32670;
    wire N__32669;
    wire N__32668;
    wire N__32667;
    wire N__32666;
    wire N__32665;
    wire N__32664;
    wire N__32663;
    wire N__32662;
    wire N__32661;
    wire N__32660;
    wire N__32659;
    wire N__32658;
    wire N__32657;
    wire N__32656;
    wire N__32655;
    wire N__32654;
    wire N__32653;
    wire N__32652;
    wire N__32649;
    wire N__32648;
    wire N__32647;
    wire N__32644;
    wire N__32635;
    wire N__32626;
    wire N__32617;
    wire N__32616;
    wire N__32613;
    wire N__32612;
    wire N__32611;
    wire N__32610;
    wire N__32609;
    wire N__32608;
    wire N__32607;
    wire N__32606;
    wire N__32605;
    wire N__32602;
    wire N__32601;
    wire N__32600;
    wire N__32599;
    wire N__32598;
    wire N__32595;
    wire N__32594;
    wire N__32591;
    wire N__32590;
    wire N__32587;
    wire N__32584;
    wire N__32581;
    wire N__32578;
    wire N__32575;
    wire N__32574;
    wire N__32573;
    wire N__32572;
    wire N__32571;
    wire N__32568;
    wire N__32559;
    wire N__32556;
    wire N__32555;
    wire N__32554;
    wire N__32553;
    wire N__32552;
    wire N__32549;
    wire N__32540;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32498;
    wire N__32497;
    wire N__32492;
    wire N__32489;
    wire N__32482;
    wire N__32475;
    wire N__32466;
    wire N__32453;
    wire N__32448;
    wire N__32443;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32419;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32399;
    wire N__32396;
    wire N__32395;
    wire N__32392;
    wire N__32389;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32377;
    wire N__32374;
    wire N__32373;
    wire N__32372;
    wire N__32369;
    wire N__32368;
    wire N__32365;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32349;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32328;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32312;
    wire N__32309;
    wire N__32308;
    wire N__32305;
    wire N__32302;
    wire N__32297;
    wire N__32296;
    wire N__32295;
    wire N__32294;
    wire N__32287;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32275;
    wire N__32272;
    wire N__32267;
    wire N__32266;
    wire N__32263;
    wire N__32262;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32231;
    wire N__32230;
    wire N__32229;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32221;
    wire N__32216;
    wire N__32213;
    wire N__32210;
    wire N__32207;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32191;
    wire N__32190;
    wire N__32189;
    wire N__32188;
    wire N__32187;
    wire N__32186;
    wire N__32185;
    wire N__32184;
    wire N__32183;
    wire N__32182;
    wire N__32181;
    wire N__32180;
    wire N__32179;
    wire N__32178;
    wire N__32177;
    wire N__32176;
    wire N__32175;
    wire N__32174;
    wire N__32173;
    wire N__32172;
    wire N__32169;
    wire N__32168;
    wire N__32167;
    wire N__32166;
    wire N__32165;
    wire N__32156;
    wire N__32147;
    wire N__32140;
    wire N__32131;
    wire N__32122;
    wire N__32119;
    wire N__32116;
    wire N__32115;
    wire N__32114;
    wire N__32113;
    wire N__32112;
    wire N__32111;
    wire N__32110;
    wire N__32109;
    wire N__32100;
    wire N__32097;
    wire N__32086;
    wire N__32083;
    wire N__32076;
    wire N__32067;
    wire N__32064;
    wire N__32059;
    wire N__32056;
    wire N__32045;
    wire N__32042;
    wire N__32041;
    wire N__32040;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32022;
    wire N__32017;
    wire N__32012;
    wire N__32009;
    wire N__32008;
    wire N__32007;
    wire N__32006;
    wire N__32005;
    wire N__32004;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31996;
    wire N__31995;
    wire N__31994;
    wire N__31993;
    wire N__31992;
    wire N__31991;
    wire N__31990;
    wire N__31989;
    wire N__31988;
    wire N__31987;
    wire N__31986;
    wire N__31985;
    wire N__31984;
    wire N__31983;
    wire N__31982;
    wire N__31981;
    wire N__31980;
    wire N__31979;
    wire N__31978;
    wire N__31977;
    wire N__31976;
    wire N__31975;
    wire N__31974;
    wire N__31973;
    wire N__31972;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31968;
    wire N__31967;
    wire N__31966;
    wire N__31965;
    wire N__31964;
    wire N__31963;
    wire N__31960;
    wire N__31959;
    wire N__31958;
    wire N__31957;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31943;
    wire N__31942;
    wire N__31941;
    wire N__31940;
    wire N__31939;
    wire N__31938;
    wire N__31937;
    wire N__31932;
    wire N__31925;
    wire N__31922;
    wire N__31913;
    wire N__31912;
    wire N__31911;
    wire N__31910;
    wire N__31909;
    wire N__31908;
    wire N__31907;
    wire N__31906;
    wire N__31905;
    wire N__31904;
    wire N__31903;
    wire N__31902;
    wire N__31901;
    wire N__31900;
    wire N__31899;
    wire N__31898;
    wire N__31895;
    wire N__31894;
    wire N__31885;
    wire N__31882;
    wire N__31865;
    wire N__31854;
    wire N__31849;
    wire N__31838;
    wire N__31835;
    wire N__31834;
    wire N__31833;
    wire N__31830;
    wire N__31823;
    wire N__31816;
    wire N__31815;
    wire N__31814;
    wire N__31813;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31801;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31781;
    wire N__31780;
    wire N__31779;
    wire N__31778;
    wire N__31777;
    wire N__31776;
    wire N__31775;
    wire N__31774;
    wire N__31773;
    wire N__31772;
    wire N__31771;
    wire N__31770;
    wire N__31769;
    wire N__31766;
    wire N__31765;
    wire N__31764;
    wire N__31761;
    wire N__31750;
    wire N__31749;
    wire N__31748;
    wire N__31747;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31731;
    wire N__31722;
    wire N__31719;
    wire N__31706;
    wire N__31701;
    wire N__31698;
    wire N__31693;
    wire N__31684;
    wire N__31679;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31656;
    wire N__31645;
    wire N__31638;
    wire N__31635;
    wire N__31630;
    wire N__31625;
    wire N__31616;
    wire N__31603;
    wire N__31584;
    wire N__31565;
    wire N__31562;
    wire N__31561;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31510;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31498;
    wire N__31493;
    wire N__31492;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31480;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31462;
    wire N__31457;
    wire N__31454;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31424;
    wire N__31421;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31413;
    wire N__31410;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31392;
    wire N__31387;
    wire N__31382;
    wire N__31381;
    wire N__31376;
    wire N__31373;
    wire N__31372;
    wire N__31371;
    wire N__31368;
    wire N__31363;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31345;
    wire N__31340;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31319;
    wire N__31316;
    wire N__31315;
    wire N__31314;
    wire N__31313;
    wire N__31312;
    wire N__31311;
    wire N__31310;
    wire N__31309;
    wire N__31308;
    wire N__31307;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31276;
    wire N__31275;
    wire N__31274;
    wire N__31271;
    wire N__31266;
    wire N__31263;
    wire N__31258;
    wire N__31253;
    wire N__31252;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31237;
    wire N__31236;
    wire N__31233;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31213;
    wire N__31208;
    wire N__31205;
    wire N__31204;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31187;
    wire N__31184;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31174;
    wire N__31173;
    wire N__31170;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31138;
    wire N__31133;
    wire N__31132;
    wire N__31129;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31121;
    wire N__31118;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31100;
    wire N__31097;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31043;
    wire N__31040;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31028;
    wire N__31025;
    wire N__31024;
    wire N__31023;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31011;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30997;
    wire N__30992;
    wire N__30991;
    wire N__30986;
    wire N__30983;
    wire N__30982;
    wire N__30981;
    wire N__30976;
    wire N__30973;
    wire N__30970;
    wire N__30965;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30957;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30941;
    wire N__30940;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30923;
    wire N__30920;
    wire N__30919;
    wire N__30916;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30895;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30862;
    wire N__30861;
    wire N__30858;
    wire N__30853;
    wire N__30848;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30827;
    wire N__30826;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30812;
    wire N__30811;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30768;
    wire N__30767;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30749;
    wire N__30746;
    wire N__30745;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30730;
    wire N__30725;
    wire N__30724;
    wire N__30721;
    wire N__30720;
    wire N__30719;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30707;
    wire N__30702;
    wire N__30695;
    wire N__30694;
    wire N__30693;
    wire N__30690;
    wire N__30685;
    wire N__30680;
    wire N__30677;
    wire N__30676;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30664;
    wire N__30663;
    wire N__30660;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30644;
    wire N__30643;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30623;
    wire N__30622;
    wire N__30619;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30595;
    wire N__30592;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30575;
    wire N__30572;
    wire N__30571;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30554;
    wire N__30551;
    wire N__30550;
    wire N__30549;
    wire N__30548;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30520;
    wire N__30519;
    wire N__30518;
    wire N__30515;
    wire N__30510;
    wire N__30507;
    wire N__30502;
    wire N__30497;
    wire N__30494;
    wire N__30493;
    wire N__30490;
    wire N__30487;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30470;
    wire N__30467;
    wire N__30466;
    wire N__30465;
    wire N__30464;
    wire N__30461;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30443;
    wire N__30440;
    wire N__30439;
    wire N__30436;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30419;
    wire N__30416;
    wire N__30415;
    wire N__30410;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30382;
    wire N__30377;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30362;
    wire N__30359;
    wire N__30358;
    wire N__30353;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30338;
    wire N__30335;
    wire N__30334;
    wire N__30333;
    wire N__30330;
    wire N__30325;
    wire N__30320;
    wire N__30317;
    wire N__30316;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30304;
    wire N__30299;
    wire N__30296;
    wire N__30295;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30278;
    wire N__30275;
    wire N__30274;
    wire N__30271;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30248;
    wire N__30245;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30233;
    wire N__30230;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30218;
    wire N__30215;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30203;
    wire N__30200;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30188;
    wire N__30185;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30173;
    wire N__30170;
    wire N__30169;
    wire N__30166;
    wire N__30161;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30139;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30124;
    wire N__30119;
    wire N__30116;
    wire N__30115;
    wire N__30110;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30082;
    wire N__30079;
    wire N__30076;
    wire N__30071;
    wire N__30068;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30056;
    wire N__30053;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30041;
    wire N__30038;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30026;
    wire N__30023;
    wire N__30022;
    wire N__30019;
    wire N__30016;
    wire N__30011;
    wire N__30008;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29996;
    wire N__29993;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29978;
    wire N__29975;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29935;
    wire N__29932;
    wire N__29929;
    wire N__29924;
    wire N__29921;
    wire N__29920;
    wire N__29919;
    wire N__29916;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29899;
    wire N__29894;
    wire N__29893;
    wire N__29890;
    wire N__29889;
    wire N__29886;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29860;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29822;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29810;
    wire N__29807;
    wire N__29806;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29789;
    wire N__29786;
    wire N__29783;
    wire N__29780;
    wire N__29779;
    wire N__29778;
    wire N__29777;
    wire N__29776;
    wire N__29775;
    wire N__29774;
    wire N__29773;
    wire N__29772;
    wire N__29771;
    wire N__29766;
    wire N__29757;
    wire N__29748;
    wire N__29745;
    wire N__29738;
    wire N__29735;
    wire N__29734;
    wire N__29731;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29714;
    wire N__29713;
    wire N__29710;
    wire N__29707;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29697;
    wire N__29696;
    wire N__29693;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29669;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29653;
    wire N__29648;
    wire N__29645;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29620;
    wire N__29619;
    wire N__29616;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29588;
    wire N__29585;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29561;
    wire N__29558;
    wire N__29557;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29540;
    wire N__29537;
    wire N__29536;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29519;
    wire N__29516;
    wire N__29515;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29498;
    wire N__29495;
    wire N__29494;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29477;
    wire N__29474;
    wire N__29473;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29456;
    wire N__29453;
    wire N__29452;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29435;
    wire N__29432;
    wire N__29429;
    wire N__29428;
    wire N__29425;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29408;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29400;
    wire N__29397;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29379;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29349;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29331;
    wire N__29326;
    wire N__29321;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29287;
    wire N__29282;
    wire N__29279;
    wire N__29278;
    wire N__29277;
    wire N__29276;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29255;
    wire N__29254;
    wire N__29253;
    wire N__29252;
    wire N__29251;
    wire N__29250;
    wire N__29249;
    wire N__29248;
    wire N__29239;
    wire N__29238;
    wire N__29237;
    wire N__29236;
    wire N__29235;
    wire N__29234;
    wire N__29233;
    wire N__29232;
    wire N__29231;
    wire N__29230;
    wire N__29229;
    wire N__29228;
    wire N__29227;
    wire N__29226;
    wire N__29225;
    wire N__29224;
    wire N__29223;
    wire N__29222;
    wire N__29221;
    wire N__29220;
    wire N__29219;
    wire N__29218;
    wire N__29217;
    wire N__29208;
    wire N__29205;
    wire N__29196;
    wire N__29191;
    wire N__29182;
    wire N__29173;
    wire N__29164;
    wire N__29155;
    wire N__29150;
    wire N__29147;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29122;
    wire N__29119;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29099;
    wire N__29096;
    wire N__29095;
    wire N__29094;
    wire N__29091;
    wire N__29088;
    wire N__29085;
    wire N__29080;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29057;
    wire N__29056;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29046;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29025;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29009;
    wire N__29008;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28984;
    wire N__28983;
    wire N__28978;
    wire N__28975;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28956;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28904;
    wire N__28903;
    wire N__28902;
    wire N__28901;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28874;
    wire N__28871;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28854;
    wire N__28851;
    wire N__28844;
    wire N__28841;
    wire N__28840;
    wire N__28839;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28823;
    wire N__28820;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28784;
    wire N__28783;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28773;
    wire N__28768;
    wire N__28763;
    wire N__28760;
    wire N__28759;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28739;
    wire N__28732;
    wire N__28729;
    wire N__28724;
    wire N__28721;
    wire N__28718;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28710;
    wire N__28709;
    wire N__28706;
    wire N__28703;
    wire N__28698;
    wire N__28695;
    wire N__28690;
    wire N__28685;
    wire N__28684;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28676;
    wire N__28675;
    wire N__28672;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28645;
    wire N__28638;
    wire N__28633;
    wire N__28630;
    wire N__28625;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28617;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28587;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28571;
    wire N__28570;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28552;
    wire N__28547;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28521;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28505;
    wire N__28504;
    wire N__28503;
    wire N__28500;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28484;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28472;
    wire N__28469;
    wire N__28466;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28436;
    wire N__28435;
    wire N__28434;
    wire N__28433;
    wire N__28430;
    wire N__28427;
    wire N__28424;
    wire N__28421;
    wire N__28418;
    wire N__28415;
    wire N__28412;
    wire N__28409;
    wire N__28404;
    wire N__28401;
    wire N__28396;
    wire N__28393;
    wire N__28388;
    wire N__28385;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28355;
    wire N__28352;
    wire N__28351;
    wire N__28350;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28334;
    wire N__28331;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28323;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28307;
    wire N__28306;
    wire N__28305;
    wire N__28302;
    wire N__28297;
    wire N__28296;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28277;
    wire N__28274;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28266;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28250;
    wire N__28249;
    wire N__28248;
    wire N__28245;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28217;
    wire N__28214;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28206;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28176;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28160;
    wire N__28157;
    wire N__28156;
    wire N__28155;
    wire N__28154;
    wire N__28151;
    wire N__28144;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28132;
    wire N__28127;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28112;
    wire N__28111;
    wire N__28108;
    wire N__28107;
    wire N__28106;
    wire N__28103;
    wire N__28100;
    wire N__28093;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28049;
    wire N__28046;
    wire N__28045;
    wire N__28044;
    wire N__28043;
    wire N__28040;
    wire N__28035;
    wire N__28032;
    wire N__28027;
    wire N__28022;
    wire N__28019;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27983;
    wire N__27982;
    wire N__27981;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27961;
    wire N__27956;
    wire N__27953;
    wire N__27952;
    wire N__27951;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27935;
    wire N__27932;
    wire N__27931;
    wire N__27926;
    wire N__27925;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27911;
    wire N__27910;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27895;
    wire N__27894;
    wire N__27889;
    wire N__27886;
    wire N__27881;
    wire N__27878;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27870;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27854;
    wire N__27851;
    wire N__27850;
    wire N__27845;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27826;
    wire N__27821;
    wire N__27818;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27796;
    wire N__27791;
    wire N__27790;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27773;
    wire N__27772;
    wire N__27769;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27752;
    wire N__27751;
    wire N__27750;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27736;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27710;
    wire N__27707;
    wire N__27704;
    wire N__27703;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27683;
    wire N__27682;
    wire N__27681;
    wire N__27678;
    wire N__27677;
    wire N__27674;
    wire N__27671;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27635;
    wire N__27632;
    wire N__27631;
    wire N__27628;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27613;
    wire N__27608;
    wire N__27607;
    wire N__27606;
    wire N__27601;
    wire N__27598;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27580;
    wire N__27575;
    wire N__27572;
    wire N__27571;
    wire N__27570;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27554;
    wire N__27551;
    wire N__27550;
    wire N__27549;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27531;
    wire N__27524;
    wire N__27521;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27513;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27481;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27469;
    wire N__27466;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27445;
    wire N__27442;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27410;
    wire N__27407;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27392;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27380;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27208;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27185;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27164;
    wire N__27161;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27098;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27080;
    wire N__27079;
    wire N__27076;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27059;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27005;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26993;
    wire N__26992;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26980;
    wire N__26977;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26960;
    wire N__26959;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26945;
    wire N__26942;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26926;
    wire N__26921;
    wire N__26918;
    wire N__26917;
    wire N__26914;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26897;
    wire N__26896;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26872;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26852;
    wire N__26851;
    wire N__26848;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26822;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26801;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26783;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26750;
    wire N__26747;
    wire N__26744;
    wire N__26741;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26723;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26675;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26657;
    wire N__26654;
    wire N__26651;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26462;
    wire N__26459;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26359;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26344;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26332;
    wire N__26331;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26308;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26209;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26197;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26185;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26170;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26147;
    wire N__26146;
    wire N__26141;
    wire N__26138;
    wire N__26137;
    wire N__26134;
    wire N__26131;
    wire N__26126;
    wire N__26123;
    wire N__26122;
    wire N__26117;
    wire N__26114;
    wire N__26111;
    wire N__26110;
    wire N__26105;
    wire N__26102;
    wire N__26101;
    wire N__26100;
    wire N__26097;
    wire N__26094;
    wire N__26091;
    wire N__26088;
    wire N__26085;
    wire N__26078;
    wire N__26077;
    wire N__26074;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26061;
    wire N__26060;
    wire N__26053;
    wire N__26050;
    wire N__26045;
    wire N__26042;
    wire N__26041;
    wire N__26038;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25987;
    wire N__25986;
    wire N__25983;
    wire N__25980;
    wire N__25975;
    wire N__25970;
    wire N__25969;
    wire N__25968;
    wire N__25965;
    wire N__25960;
    wire N__25955;
    wire N__25954;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25931;
    wire N__25928;
    wire N__25927;
    wire N__25926;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25914;
    wire N__25907;
    wire N__25904;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25889;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25877;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25862;
    wire N__25859;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25846;
    wire N__25841;
    wire N__25838;
    wire N__25837;
    wire N__25836;
    wire N__25833;
    wire N__25828;
    wire N__25823;
    wire N__25822;
    wire N__25821;
    wire N__25818;
    wire N__25813;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25735;
    wire N__25734;
    wire N__25733;
    wire N__25732;
    wire N__25721;
    wire N__25720;
    wire N__25719;
    wire N__25718;
    wire N__25717;
    wire N__25716;
    wire N__25713;
    wire N__25702;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25690;
    wire N__25689;
    wire N__25688;
    wire N__25687;
    wire N__25686;
    wire N__25685;
    wire N__25684;
    wire N__25683;
    wire N__25682;
    wire N__25671;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25601;
    wire N__25598;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25571;
    wire N__25568;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25546;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25510;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25498;
    wire N__25497;
    wire N__25496;
    wire N__25495;
    wire N__25494;
    wire N__25493;
    wire N__25492;
    wire N__25491;
    wire N__25490;
    wire N__25489;
    wire N__25488;
    wire N__25487;
    wire N__25486;
    wire N__25485;
    wire N__25484;
    wire N__25483;
    wire N__25480;
    wire N__25463;
    wire N__25446;
    wire N__25443;
    wire N__25442;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25412;
    wire N__25409;
    wire N__25406;
    wire N__25403;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25372;
    wire N__25369;
    wire N__25366;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25345;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25328;
    wire N__25325;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25298;
    wire N__25295;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25273;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25106;
    wire N__25105;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25093;
    wire N__25092;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25076;
    wire N__25075;
    wire N__25072;
    wire N__25071;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25030;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__24998;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24938;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24890;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24854;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24656;
    wire N__24653;
    wire N__24650;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24554;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24541;
    wire N__24540;
    wire N__24539;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24514;
    wire N__24513;
    wire N__24512;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24439;
    wire N__24436;
    wire N__24433;
    wire N__24430;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24403;
    wire N__24402;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24379;
    wire N__24374;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24346;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24331;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24316;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24296;
    wire N__24293;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24218;
    wire N__24215;
    wire N__24212;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24131;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24080;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24056;
    wire N__24055;
    wire N__24054;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24031;
    wire N__24030;
    wire N__24027;
    wire N__24020;
    wire N__24019;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24011;
    wire N__24010;
    wire N__24009;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23986;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23942;
    wire N__23941;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23917;
    wire N__23916;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23904;
    wire N__23903;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23836;
    wire N__23831;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23818;
    wire N__23817;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23791;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23768;
    wire N__23765;
    wire N__23762;
    wire N__23759;
    wire N__23758;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23731;
    wire N__23728;
    wire N__23725;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23710;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23569;
    wire N__23566;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23550;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23513;
    wire N__23510;
    wire N__23509;
    wire N__23506;
    wire N__23505;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23420;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23287;
    wire N__23284;
    wire N__23283;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23271;
    wire N__23268;
    wire N__23261;
    wire N__23260;
    wire N__23259;
    wire N__23258;
    wire N__23257;
    wire N__23256;
    wire N__23255;
    wire N__23254;
    wire N__23253;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23235;
    wire N__23234;
    wire N__23233;
    wire N__23232;
    wire N__23231;
    wire N__23230;
    wire N__23229;
    wire N__23228;
    wire N__23227;
    wire N__23224;
    wire N__23223;
    wire N__23222;
    wire N__23217;
    wire N__23212;
    wire N__23207;
    wire N__23204;
    wire N__23193;
    wire N__23190;
    wire N__23189;
    wire N__23188;
    wire N__23187;
    wire N__23186;
    wire N__23185;
    wire N__23184;
    wire N__23183;
    wire N__23182;
    wire N__23181;
    wire N__23168;
    wire N__23165;
    wire N__23160;
    wire N__23159;
    wire N__23156;
    wire N__23149;
    wire N__23144;
    wire N__23141;
    wire N__23128;
    wire N__23123;
    wire N__23120;
    wire N__23117;
    wire N__23114;
    wire N__23111;
    wire N__23106;
    wire N__23103;
    wire N__23084;
    wire N__23083;
    wire N__23082;
    wire N__23081;
    wire N__23078;
    wire N__23077;
    wire N__23076;
    wire N__23075;
    wire N__23074;
    wire N__23073;
    wire N__23068;
    wire N__23065;
    wire N__23064;
    wire N__23063;
    wire N__23058;
    wire N__23055;
    wire N__23054;
    wire N__23053;
    wire N__23052;
    wire N__23051;
    wire N__23050;
    wire N__23049;
    wire N__23048;
    wire N__23047;
    wire N__23046;
    wire N__23045;
    wire N__23044;
    wire N__23043;
    wire N__23042;
    wire N__23041;
    wire N__23040;
    wire N__23039;
    wire N__23038;
    wire N__23037;
    wire N__23036;
    wire N__23035;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23021;
    wire N__23016;
    wire N__23011;
    wire N__23002;
    wire N__22997;
    wire N__22990;
    wire N__22977;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22955;
    wire N__22950;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22913;
    wire N__22912;
    wire N__22909;
    wire N__22908;
    wire N__22905;
    wire N__22904;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22883;
    wire N__22874;
    wire N__22873;
    wire N__22870;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22862;
    wire N__22859;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22832;
    wire N__22831;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22800;
    wire N__22793;
    wire N__22792;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22766;
    wire N__22763;
    wire N__22758;
    wire N__22755;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22732;
    wire N__22731;
    wire N__22728;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22718;
    wire N__22715;
    wire N__22710;
    wire N__22703;
    wire N__22700;
    wire N__22699;
    wire N__22696;
    wire N__22695;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22633;
    wire N__22632;
    wire N__22631;
    wire N__22630;
    wire N__22629;
    wire N__22628;
    wire N__22627;
    wire N__22626;
    wire N__22625;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22617;
    wire N__22616;
    wire N__22615;
    wire N__22614;
    wire N__22613;
    wire N__22612;
    wire N__22611;
    wire N__22610;
    wire N__22609;
    wire N__22608;
    wire N__22607;
    wire N__22606;
    wire N__22603;
    wire N__22602;
    wire N__22599;
    wire N__22598;
    wire N__22597;
    wire N__22582;
    wire N__22577;
    wire N__22566;
    wire N__22565;
    wire N__22564;
    wire N__22561;
    wire N__22556;
    wire N__22553;
    wire N__22552;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22541;
    wire N__22538;
    wire N__22533;
    wire N__22528;
    wire N__22525;
    wire N__22520;
    wire N__22515;
    wire N__22510;
    wire N__22507;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22472;
    wire N__22465;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22435;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22400;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22385;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22367;
    wire N__22364;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22048;
    wire N__22047;
    wire N__22046;
    wire N__22045;
    wire N__22044;
    wire N__22043;
    wire N__22042;
    wire N__22041;
    wire N__22038;
    wire N__22037;
    wire N__22034;
    wire N__22033;
    wire N__22030;
    wire N__22029;
    wire N__22026;
    wire N__22025;
    wire N__22022;
    wire N__22021;
    wire N__22018;
    wire N__22017;
    wire N__22014;
    wire N__22013;
    wire N__22012;
    wire N__22009;
    wire N__22008;
    wire N__21993;
    wire N__21976;
    wire N__21969;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21598;
    wire N__21597;
    wire N__21596;
    wire N__21593;
    wire N__21590;
    wire N__21587;
    wire N__21584;
    wire N__21575;
    wire N__21574;
    wire N__21571;
    wire N__21570;
    wire N__21567;
    wire N__21566;
    wire N__21563;
    wire N__21560;
    wire N__21557;
    wire N__21554;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21517;
    wire N__21516;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21504;
    wire N__21497;
    wire N__21494;
    wire N__21493;
    wire N__21492;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21480;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21466;
    wire N__21463;
    wire N__21462;
    wire N__21459;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21447;
    wire N__21440;
    wire N__21439;
    wire N__21436;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21409;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21397;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21389;
    wire N__21386;
    wire N__21381;
    wire N__21378;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21364;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21356;
    wire N__21353;
    wire N__21348;
    wire N__21345;
    wire N__21338;
    wire N__21335;
    wire N__21334;
    wire N__21333;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21321;
    wire N__21314;
    wire N__21313;
    wire N__21310;
    wire N__21309;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21296;
    wire N__21293;
    wire N__21288;
    wire N__21285;
    wire N__21280;
    wire N__21277;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21244;
    wire N__21241;
    wire N__21240;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21228;
    wire N__21225;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21187;
    wire N__21186;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21174;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21157;
    wire N__21156;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21144;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21130;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21119;
    wire N__21116;
    wire N__21111;
    wire N__21108;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21091;
    wire N__21090;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21061;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21048;
    wire N__21041;
    wire N__21038;
    wire N__21037;
    wire N__21036;
    wire N__21033;
    wire N__21032;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21011;
    wire N__21010;
    wire N__21009;
    wire N__21006;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20988;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20974;
    wire N__20973;
    wire N__20972;
    wire N__20969;
    wire N__20966;
    wire N__20961;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20947;
    wire N__20946;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20936;
    wire N__20933;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20884;
    wire N__20881;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20846;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20838;
    wire N__20835;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20791;
    wire N__20788;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20704;
    wire N__20701;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20669;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20650;
    wire N__20645;
    wire N__20642;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20617;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20582;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20567;
    wire N__20564;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20552;
    wire N__20549;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20524;
    wire N__20521;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20503;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20467;
    wire N__20462;
    wire N__20461;
    wire N__20458;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20429;
    wire N__20426;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20401;
    wire N__20396;
    wire N__20393;
    wire N__20390;
    wire N__20387;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20339;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20309;
    wire N__20308;
    wire N__20305;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20290;
    wire N__20285;
    wire N__20282;
    wire N__20281;
    wire N__20278;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20251;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20237;
    wire N__20234;
    wire N__20233;
    wire N__20230;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20218;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20206;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20194;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20182;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20159;
    wire N__20156;
    wire N__20155;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20099;
    wire N__20096;
    wire N__20095;
    wire N__20090;
    wire N__20087;
    wire N__20084;
    wire N__20083;
    wire N__20078;
    wire N__20075;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20036;
    wire N__20033;
    wire N__20032;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19904;
    wire N__19901;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19822;
    wire N__19819;
    wire N__19818;
    wire N__19815;
    wire N__19810;
    wire N__19809;
    wire N__19808;
    wire N__19807;
    wire N__19804;
    wire N__19803;
    wire N__19800;
    wire N__19799;
    wire N__19798;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19769;
    wire N__19760;
    wire N__19757;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19745;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19737;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19718;
    wire N__19715;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19700;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19685;
    wire N__19682;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19654;
    wire N__19653;
    wire N__19650;
    wire N__19645;
    wire N__19642;
    wire N__19637;
    wire N__19636;
    wire N__19635;
    wire N__19632;
    wire N__19627;
    wire N__19624;
    wire N__19619;
    wire N__19618;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19595;
    wire N__19594;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19510;
    wire N__19509;
    wire N__19504;
    wire N__19501;
    wire N__19496;
    wire N__19495;
    wire N__19494;
    wire N__19491;
    wire N__19490;
    wire N__19489;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19475;
    wire N__19472;
    wire N__19465;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19448;
    wire N__19447;
    wire N__19446;
    wire N__19445;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18881;
    wire N__18878;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18848;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18730;
    wire N__18729;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18661;
    wire N__18660;
    wire N__18659;
    wire N__18658;
    wire N__18657;
    wire N__18656;
    wire N__18655;
    wire N__18654;
    wire N__18653;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18621;
    wire N__18618;
    wire N__18609;
    wire N__18606;
    wire N__18599;
    wire N__18592;
    wire N__18585;
    wire N__18580;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire GNDG0;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire bfn_1_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire bfn_1_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire N_42_i_i;
    wire un7_start_stop_0_a2;
    wire bfn_2_13_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire bfn_2_14_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire bfn_2_15_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire bfn_2_16_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.N_159 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.N_96_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_0_3 ;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_7;
    wire pwm_duty_input_6;
    wire pwm_duty_input_8;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire bfn_3_17_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire bfn_3_18_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire bfn_3_19_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire bfn_3_20_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.N_98 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire pwm_duty_input_3;
    wire pwm_duty_input_4;
    wire pwm_duty_input_5;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ;
    wire bfn_3_24_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire bfn_3_25_0_;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire bfn_3_26_0_;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.N_77_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire bfn_4_23_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ;
    wire bfn_4_24_0_;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire bfn_4_25_0_;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_ ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16_cascade_ ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.N_44_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.N_46 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_5_25_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_5_26_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire bfn_5_27_0_;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire bfn_7_23_0_;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire bfn_7_24_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire il_max_comp1_c;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ;
    wire bfn_8_5_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_8_6_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_8_7_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_8_8_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_8_9_0_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_8_10_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire bfn_8_11_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire elapsed_time_ns_1_RNI58DN9_0_27_cascade_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.N_16 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire elapsed_time_ns_1_RNI24CN9_0_15_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire elapsed_time_ns_1_RNITUBN9_0_10_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire bfn_9_15_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_9_16_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_9_17_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_9_18_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \current_shift_inst.control_input_18 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_9_20_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \pwm_generator_inst.threshold_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_9_24_0_;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_9_25_0_;
    wire \pwm_generator_inst.threshold_9 ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire s3_phy_c;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_10_7_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_10_8_0_;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire bfn_10_9_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt26 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire bfn_10_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire bfn_10_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire bfn_10_14_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire bfn_10_15_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.N_202_i ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire \delay_measurement_inst.delay_hc_timer.N_203_i ;
    wire il_max_comp1_D1;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.N_1304_i ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire bfn_10_24_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_10_25_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_df30_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire bfn_11_8_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire bfn_11_9_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire bfn_11_10_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_11_11_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire start_stop_c;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire \phase_controller_inst2.start_timer_tr_RNO_0_0 ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.start_timer_hc_0_sqmuxa ;
    wire \phase_controller_inst2.state_RNIG7JFZ0Z_2 ;
    wire il_min_comp2_c;
    wire il_max_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt28 ;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire elapsed_time_ns_1_RNI7ADN9_0_29_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.un1_start_g ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire bfn_12_15_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire bfn_12_16_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_12_17_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire bfn_12_18_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire il_min_comp1_c;
    wire il_min_comp1_D1;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire s4_phy_c;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire delay_hc_input_c_g;
    wire \pll_inst.red_c_i ;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.state_RNI9M3OZ0Z_0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst2.stoper_tr.un4_running_df30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13_cascade_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ;
    wire bfn_13_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_13_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_13_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_13_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.N_205_i ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire state_ns_i_a2_1;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.start_timer_hc_0_sqmuxa ;
    wire il_max_comp1_D2;
    wire \current_shift_inst.timer_s1.N_162_i ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ;
    wire bfn_14_8_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire bfn_14_9_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_14_10_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_14_11_0_;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire elapsed_time_ns_1_RNIVAQBB_0_30_cascade_;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire elapsed_time_ns_1_RNI0CQBB_0_31_cascade_;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire bfn_14_13_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire bfn_14_14_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire phase_controller_inst1_state_4;
    wire \phase_controller_inst1.time_passed_RNIE87F ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire il_min_comp1_D2;
    wire \phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire s1_phy_c;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire s2_phy_c;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_15_7_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_15_8_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire bfn_15_9_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_15_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_15_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_15_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_15_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_204_i ;
    wire \current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire bfn_15_18_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire bfn_15_19_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire bfn_15_20_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire bfn_15_21_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire T12_c;
    wire T45_c;
    wire state_3;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire T01_c;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire T23_c;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire elapsed_time_ns_1_RNIU7OBB_0_11_cascade_;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire elapsed_time_ns_1_RNIT6OBB_0_10_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_16_11_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_16_12_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire bfn_16_13_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire bfn_16_14_0_;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire bfn_16_15_0_;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_16_16_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_16_17_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.time_passed_RNI7NN7 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire elapsed_time_ns_1_RNIV9PBB_0_21_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire elapsed_time_ns_1_RNI0BPBB_0_22_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_17_10_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_17_11_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_17_12_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire bfn_17_13_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_17_19_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_17_20_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_17_21_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_163_i ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire \phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_df30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ;
    wire \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire elapsed_time_ns_1_RNI5FOBB_0_18_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire bfn_18_14_0_;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire bfn_18_15_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire bfn_18_16_0_;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire bfn_18_17_0_;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.N_162_i_g ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.un1_start_g ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire clk_100mhz_0;
    wire \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ;
    wire red_c_g;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire N_19_1;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire _gnd_net_;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__30875),
            .RESETB(N__32915),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37930),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37905),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__25490,N__25498,N__25489,N__25496,N__25488,N__25495,N__25487,N__25497,N__25484,N__25491,N__25483,N__25492,N__25486,N__25493,N__25485,N__25494}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__37929,dangling_wire_45,N__37928}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37904),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37897),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__46183,N__46176,N__46181,N__46175,N__46182,N__46174,N__46184,N__46171,N__46177,N__46170,N__46178,N__46172,N__46179,N__46173,N__46180}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,N__37903,N__37900,dangling_wire_102,dangling_wire_103,dangling_wire_104,N__37898,N__37902,N__37899,N__37901}),
            .OHOLDTOP(),
            .O({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37980),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37823),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .ADDSUBBOT(),
            .A({dangling_wire_136,N__46231,N__46234,N__46232,N__46235,N__46233,N__19655,N__19593,N__19637,N__19618,N__20281,N__20309,N__20338,N__19685,N__19700,N__19718}),
            .C({dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}),
            .B({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,N__37829,N__37826,dangling_wire_160,dangling_wire_161,dangling_wire_162,N__37824,N__37828,N__37825,N__37827}),
            .OHOLDTOP(),
            .O({dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__37979),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__37976),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .ADDSUBBOT(),
            .A({dangling_wire_185,N__25499,N__25538,N__25568,N__25598,N__25631,N__25136,N__25166,N__25199,N__25232,N__25265,N__25295,N__25325,N__25355,N__25384,N__24998}),
            .C({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .B({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__37978,dangling_wire_215,N__37977}),
            .OHOLDTOP(),
            .O({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__48450),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__48452),
            .DIN(N__48451),
            .DOUT(N__48450),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__48452),
            .PADOUT(N__48451),
            .PADIN(N__48450),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T01_obuf_iopad (
            .OE(N__48441),
            .DIN(N__48440),
            .DOUT(N__48439),
            .PACKAGEPIN(T01));
    defparam T01_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T01_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T01_obuf_preio (
            .PADOEN(N__48441),
            .PADOUT(N__48440),
            .PADIN(N__48439),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36608),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__48432),
            .DIN(N__48431),
            .DOUT(N__48430),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__48432),
            .PADOUT(N__48431),
            .PADIN(N__48430),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__48423),
            .DIN(N__48422),
            .DOUT(N__48421),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__48423),
            .PADOUT(N__48422),
            .PADIN(N__48421),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T23_obuf_iopad (
            .OE(N__48414),
            .DIN(N__48413),
            .DOUT(N__48412),
            .PACKAGEPIN(T23));
    defparam T23_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T23_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T23_obuf_preio (
            .PADOEN(N__48414),
            .PADOUT(N__48413),
            .PADIN(N__48412),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36545),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__48405),
            .DIN(N__48404),
            .DOUT(N__48403),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__48405),
            .PADOUT(N__48404),
            .PADIN(N__48403),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26735),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__48396),
            .DIN(N__48395),
            .DOUT(N__48394),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__48396),
            .PADOUT(N__48395),
            .PADIN(N__48394),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__48387),
            .DIN(N__48386),
            .DOUT(N__48385),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__48387),
            .PADOUT(N__48386),
            .PADIN(N__48385),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34814),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T12_obuf_iopad (
            .OE(N__48378),
            .DIN(N__48377),
            .DOUT(N__48376),
            .PACKAGEPIN(T12));
    defparam T12_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T12_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T12_obuf_preio (
            .PADOEN(N__48378),
            .PADOUT(N__48377),
            .PADIN(N__48376),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36749),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__48369),
            .DIN(N__48368),
            .DOUT(N__48367),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__48369),
            .PADOUT(N__48368),
            .PADIN(N__48367),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__48360),
            .DIN(N__48359),
            .DOUT(N__48358),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__48360),
            .PADOUT(N__48359),
            .PADIN(N__48358),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__34871),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__48351),
            .DIN(N__48350),
            .DOUT(N__48349),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__48351),
            .PADOUT(N__48350),
            .PADIN(N__48349),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__32978),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__48342),
            .DIN(N__48341),
            .DOUT(N__48340),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__48342),
            .PADOUT(N__48341),
            .PADIN(N__48340),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__48333),
            .DIN(N__48332),
            .DOUT(N__48331),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__48333),
            .PADOUT(N__48332),
            .PADIN(N__48331),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__26714),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD T45_obuf_iopad (
            .OE(N__48324),
            .DIN(N__48323),
            .DOUT(N__48322),
            .PACKAGEPIN(T45));
    defparam T45_obuf_preio.NEG_TRIGGER=1'b0;
    defparam T45_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO T45_obuf_preio (
            .PADOEN(N__48324),
            .PADOUT(N__48323),
            .PADIN(N__48322),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__36728),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__48315),
            .DIN(N__48314),
            .DOUT(N__48313),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__48315),
            .PADOUT(N__48314),
            .PADIN(N__48313),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__48306),
            .DIN(N__48305),
            .DOUT(N__48304),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__48306),
            .PADOUT(N__48305),
            .PADIN(N__48304),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__11505 (
            .O(N__48287),
            .I(N__48281));
    InMux I__11504 (
            .O(N__48286),
            .I(N__48278));
    InMux I__11503 (
            .O(N__48285),
            .I(N__48275));
    InMux I__11502 (
            .O(N__48284),
            .I(N__48272));
    LocalMux I__11501 (
            .O(N__48281),
            .I(N__48269));
    LocalMux I__11500 (
            .O(N__48278),
            .I(N__48266));
    LocalMux I__11499 (
            .O(N__48275),
            .I(N__48263));
    LocalMux I__11498 (
            .O(N__48272),
            .I(N__48260));
    Span4Mux_v I__11497 (
            .O(N__48269),
            .I(N__48257));
    Span4Mux_h I__11496 (
            .O(N__48266),
            .I(N__48254));
    Span4Mux_h I__11495 (
            .O(N__48263),
            .I(N__48251));
    Span4Mux_h I__11494 (
            .O(N__48260),
            .I(N__48248));
    Span4Mux_h I__11493 (
            .O(N__48257),
            .I(N__48245));
    Span4Mux_h I__11492 (
            .O(N__48254),
            .I(N__48242));
    Span4Mux_h I__11491 (
            .O(N__48251),
            .I(N__48239));
    Span4Mux_v I__11490 (
            .O(N__48248),
            .I(N__48236));
    Odrv4 I__11489 (
            .O(N__48245),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__11488 (
            .O(N__48242),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__11487 (
            .O(N__48239),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__11486 (
            .O(N__48236),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__11485 (
            .O(N__48227),
            .I(N__48223));
    InMux I__11484 (
            .O(N__48226),
            .I(N__48219));
    LocalMux I__11483 (
            .O(N__48223),
            .I(N__48216));
    InMux I__11482 (
            .O(N__48222),
            .I(N__48213));
    LocalMux I__11481 (
            .O(N__48219),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    Odrv4 I__11480 (
            .O(N__48216),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    LocalMux I__11479 (
            .O(N__48213),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    CascadeMux I__11478 (
            .O(N__48206),
            .I(N__48190));
    CascadeMux I__11477 (
            .O(N__48205),
            .I(N__48173));
    CascadeMux I__11476 (
            .O(N__48204),
            .I(N__48170));
    InMux I__11475 (
            .O(N__48203),
            .I(N__48160));
    InMux I__11474 (
            .O(N__48202),
            .I(N__48160));
    InMux I__11473 (
            .O(N__48201),
            .I(N__48160));
    InMux I__11472 (
            .O(N__48200),
            .I(N__48160));
    InMux I__11471 (
            .O(N__48199),
            .I(N__48155));
    InMux I__11470 (
            .O(N__48198),
            .I(N__48155));
    InMux I__11469 (
            .O(N__48197),
            .I(N__48133));
    InMux I__11468 (
            .O(N__48196),
            .I(N__48133));
    InMux I__11467 (
            .O(N__48195),
            .I(N__48133));
    InMux I__11466 (
            .O(N__48194),
            .I(N__48133));
    InMux I__11465 (
            .O(N__48193),
            .I(N__48133));
    InMux I__11464 (
            .O(N__48190),
            .I(N__48118));
    InMux I__11463 (
            .O(N__48189),
            .I(N__48118));
    InMux I__11462 (
            .O(N__48188),
            .I(N__48118));
    InMux I__11461 (
            .O(N__48187),
            .I(N__48118));
    InMux I__11460 (
            .O(N__48186),
            .I(N__48118));
    InMux I__11459 (
            .O(N__48185),
            .I(N__48105));
    InMux I__11458 (
            .O(N__48184),
            .I(N__48105));
    InMux I__11457 (
            .O(N__48183),
            .I(N__48105));
    InMux I__11456 (
            .O(N__48182),
            .I(N__48105));
    InMux I__11455 (
            .O(N__48181),
            .I(N__48105));
    InMux I__11454 (
            .O(N__48180),
            .I(N__48102));
    CascadeMux I__11453 (
            .O(N__48179),
            .I(N__48092));
    InMux I__11452 (
            .O(N__48178),
            .I(N__48080));
    InMux I__11451 (
            .O(N__48177),
            .I(N__48080));
    InMux I__11450 (
            .O(N__48176),
            .I(N__48080));
    InMux I__11449 (
            .O(N__48173),
            .I(N__48073));
    InMux I__11448 (
            .O(N__48170),
            .I(N__48073));
    InMux I__11447 (
            .O(N__48169),
            .I(N__48073));
    LocalMux I__11446 (
            .O(N__48160),
            .I(N__48068));
    LocalMux I__11445 (
            .O(N__48155),
            .I(N__48068));
    InMux I__11444 (
            .O(N__48154),
            .I(N__48063));
    InMux I__11443 (
            .O(N__48153),
            .I(N__48063));
    InMux I__11442 (
            .O(N__48152),
            .I(N__48060));
    InMux I__11441 (
            .O(N__48151),
            .I(N__48057));
    InMux I__11440 (
            .O(N__48150),
            .I(N__48052));
    InMux I__11439 (
            .O(N__48149),
            .I(N__48052));
    InMux I__11438 (
            .O(N__48148),
            .I(N__48042));
    InMux I__11437 (
            .O(N__48147),
            .I(N__48042));
    InMux I__11436 (
            .O(N__48146),
            .I(N__48042));
    InMux I__11435 (
            .O(N__48145),
            .I(N__48042));
    InMux I__11434 (
            .O(N__48144),
            .I(N__48039));
    LocalMux I__11433 (
            .O(N__48133),
            .I(N__48036));
    InMux I__11432 (
            .O(N__48132),
            .I(N__48027));
    InMux I__11431 (
            .O(N__48131),
            .I(N__48027));
    InMux I__11430 (
            .O(N__48130),
            .I(N__48027));
    InMux I__11429 (
            .O(N__48129),
            .I(N__48027));
    LocalMux I__11428 (
            .O(N__48118),
            .I(N__48016));
    InMux I__11427 (
            .O(N__48117),
            .I(N__48011));
    InMux I__11426 (
            .O(N__48116),
            .I(N__48011));
    LocalMux I__11425 (
            .O(N__48105),
            .I(N__47992));
    LocalMux I__11424 (
            .O(N__48102),
            .I(N__47989));
    InMux I__11423 (
            .O(N__48101),
            .I(N__47971));
    InMux I__11422 (
            .O(N__48100),
            .I(N__47971));
    InMux I__11421 (
            .O(N__48099),
            .I(N__47971));
    InMux I__11420 (
            .O(N__48098),
            .I(N__47971));
    InMux I__11419 (
            .O(N__48097),
            .I(N__47960));
    InMux I__11418 (
            .O(N__48096),
            .I(N__47960));
    InMux I__11417 (
            .O(N__48095),
            .I(N__47960));
    InMux I__11416 (
            .O(N__48092),
            .I(N__47960));
    InMux I__11415 (
            .O(N__48091),
            .I(N__47960));
    InMux I__11414 (
            .O(N__48090),
            .I(N__47951));
    InMux I__11413 (
            .O(N__48089),
            .I(N__47951));
    InMux I__11412 (
            .O(N__48088),
            .I(N__47951));
    InMux I__11411 (
            .O(N__48087),
            .I(N__47951));
    LocalMux I__11410 (
            .O(N__48080),
            .I(N__47936));
    LocalMux I__11409 (
            .O(N__48073),
            .I(N__47936));
    Span4Mux_v I__11408 (
            .O(N__48068),
            .I(N__47936));
    LocalMux I__11407 (
            .O(N__48063),
            .I(N__47936));
    LocalMux I__11406 (
            .O(N__48060),
            .I(N__47936));
    LocalMux I__11405 (
            .O(N__48057),
            .I(N__47936));
    LocalMux I__11404 (
            .O(N__48052),
            .I(N__47936));
    InMux I__11403 (
            .O(N__48051),
            .I(N__47933));
    LocalMux I__11402 (
            .O(N__48042),
            .I(N__47928));
    LocalMux I__11401 (
            .O(N__48039),
            .I(N__47928));
    Span4Mux_v I__11400 (
            .O(N__48036),
            .I(N__47925));
    LocalMux I__11399 (
            .O(N__48027),
            .I(N__47922));
    InMux I__11398 (
            .O(N__48026),
            .I(N__47917));
    InMux I__11397 (
            .O(N__48025),
            .I(N__47917));
    InMux I__11396 (
            .O(N__48024),
            .I(N__47910));
    InMux I__11395 (
            .O(N__48023),
            .I(N__47910));
    InMux I__11394 (
            .O(N__48022),
            .I(N__47910));
    InMux I__11393 (
            .O(N__48021),
            .I(N__47903));
    InMux I__11392 (
            .O(N__48020),
            .I(N__47903));
    InMux I__11391 (
            .O(N__48019),
            .I(N__47903));
    Span4Mux_v I__11390 (
            .O(N__48016),
            .I(N__47898));
    LocalMux I__11389 (
            .O(N__48011),
            .I(N__47898));
    InMux I__11388 (
            .O(N__48010),
            .I(N__47895));
    InMux I__11387 (
            .O(N__48009),
            .I(N__47886));
    InMux I__11386 (
            .O(N__48008),
            .I(N__47886));
    InMux I__11385 (
            .O(N__48007),
            .I(N__47886));
    InMux I__11384 (
            .O(N__48006),
            .I(N__47886));
    InMux I__11383 (
            .O(N__48005),
            .I(N__47879));
    InMux I__11382 (
            .O(N__48004),
            .I(N__47879));
    InMux I__11381 (
            .O(N__48003),
            .I(N__47879));
    InMux I__11380 (
            .O(N__48002),
            .I(N__47870));
    InMux I__11379 (
            .O(N__48001),
            .I(N__47870));
    InMux I__11378 (
            .O(N__48000),
            .I(N__47870));
    InMux I__11377 (
            .O(N__47999),
            .I(N__47870));
    InMux I__11376 (
            .O(N__47998),
            .I(N__47861));
    InMux I__11375 (
            .O(N__47997),
            .I(N__47861));
    InMux I__11374 (
            .O(N__47996),
            .I(N__47861));
    InMux I__11373 (
            .O(N__47995),
            .I(N__47861));
    Span4Mux_h I__11372 (
            .O(N__47992),
            .I(N__47856));
    Span4Mux_v I__11371 (
            .O(N__47989),
            .I(N__47856));
    InMux I__11370 (
            .O(N__47988),
            .I(N__47853));
    InMux I__11369 (
            .O(N__47987),
            .I(N__47848));
    InMux I__11368 (
            .O(N__47986),
            .I(N__47848));
    InMux I__11367 (
            .O(N__47985),
            .I(N__47839));
    InMux I__11366 (
            .O(N__47984),
            .I(N__47839));
    InMux I__11365 (
            .O(N__47983),
            .I(N__47839));
    InMux I__11364 (
            .O(N__47982),
            .I(N__47839));
    InMux I__11363 (
            .O(N__47981),
            .I(N__47834));
    InMux I__11362 (
            .O(N__47980),
            .I(N__47834));
    LocalMux I__11361 (
            .O(N__47971),
            .I(N__47827));
    LocalMux I__11360 (
            .O(N__47960),
            .I(N__47827));
    LocalMux I__11359 (
            .O(N__47951),
            .I(N__47827));
    Span4Mux_v I__11358 (
            .O(N__47936),
            .I(N__47824));
    LocalMux I__11357 (
            .O(N__47933),
            .I(N__47813));
    Span4Mux_h I__11356 (
            .O(N__47928),
            .I(N__47813));
    Span4Mux_h I__11355 (
            .O(N__47925),
            .I(N__47813));
    Span4Mux_v I__11354 (
            .O(N__47922),
            .I(N__47813));
    LocalMux I__11353 (
            .O(N__47917),
            .I(N__47813));
    LocalMux I__11352 (
            .O(N__47910),
            .I(N__47806));
    LocalMux I__11351 (
            .O(N__47903),
            .I(N__47806));
    Span4Mux_h I__11350 (
            .O(N__47898),
            .I(N__47806));
    LocalMux I__11349 (
            .O(N__47895),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11348 (
            .O(N__47886),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11347 (
            .O(N__47879),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11346 (
            .O(N__47870),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11345 (
            .O(N__47861),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11344 (
            .O(N__47856),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11343 (
            .O(N__47853),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11342 (
            .O(N__47848),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11341 (
            .O(N__47839),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__11340 (
            .O(N__47834),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11339 (
            .O(N__47827),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11338 (
            .O(N__47824),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11337 (
            .O(N__47813),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__11336 (
            .O(N__47806),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    CascadeMux I__11335 (
            .O(N__47777),
            .I(N__47772));
    InMux I__11334 (
            .O(N__47776),
            .I(N__47769));
    InMux I__11333 (
            .O(N__47775),
            .I(N__47766));
    InMux I__11332 (
            .O(N__47772),
            .I(N__47763));
    LocalMux I__11331 (
            .O(N__47769),
            .I(N__47759));
    LocalMux I__11330 (
            .O(N__47766),
            .I(N__47756));
    LocalMux I__11329 (
            .O(N__47763),
            .I(N__47753));
    InMux I__11328 (
            .O(N__47762),
            .I(N__47750));
    Span4Mux_h I__11327 (
            .O(N__47759),
            .I(N__47747));
    Span4Mux_h I__11326 (
            .O(N__47756),
            .I(N__47744));
    Span4Mux_h I__11325 (
            .O(N__47753),
            .I(N__47741));
    LocalMux I__11324 (
            .O(N__47750),
            .I(N__47738));
    Span4Mux_h I__11323 (
            .O(N__47747),
            .I(N__47735));
    Span4Mux_h I__11322 (
            .O(N__47744),
            .I(N__47730));
    Span4Mux_v I__11321 (
            .O(N__47741),
            .I(N__47730));
    Odrv12 I__11320 (
            .O(N__47738),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__11319 (
            .O(N__47735),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__11318 (
            .O(N__47730),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__11317 (
            .O(N__47723),
            .I(N__47719));
    InMux I__11316 (
            .O(N__47722),
            .I(N__47715));
    LocalMux I__11315 (
            .O(N__47719),
            .I(N__47712));
    InMux I__11314 (
            .O(N__47718),
            .I(N__47709));
    LocalMux I__11313 (
            .O(N__47715),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    Odrv4 I__11312 (
            .O(N__47712),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    LocalMux I__11311 (
            .O(N__47709),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    ClkMux I__11310 (
            .O(N__47702),
            .I(N__47240));
    ClkMux I__11309 (
            .O(N__47701),
            .I(N__47240));
    ClkMux I__11308 (
            .O(N__47700),
            .I(N__47240));
    ClkMux I__11307 (
            .O(N__47699),
            .I(N__47240));
    ClkMux I__11306 (
            .O(N__47698),
            .I(N__47240));
    ClkMux I__11305 (
            .O(N__47697),
            .I(N__47240));
    ClkMux I__11304 (
            .O(N__47696),
            .I(N__47240));
    ClkMux I__11303 (
            .O(N__47695),
            .I(N__47240));
    ClkMux I__11302 (
            .O(N__47694),
            .I(N__47240));
    ClkMux I__11301 (
            .O(N__47693),
            .I(N__47240));
    ClkMux I__11300 (
            .O(N__47692),
            .I(N__47240));
    ClkMux I__11299 (
            .O(N__47691),
            .I(N__47240));
    ClkMux I__11298 (
            .O(N__47690),
            .I(N__47240));
    ClkMux I__11297 (
            .O(N__47689),
            .I(N__47240));
    ClkMux I__11296 (
            .O(N__47688),
            .I(N__47240));
    ClkMux I__11295 (
            .O(N__47687),
            .I(N__47240));
    ClkMux I__11294 (
            .O(N__47686),
            .I(N__47240));
    ClkMux I__11293 (
            .O(N__47685),
            .I(N__47240));
    ClkMux I__11292 (
            .O(N__47684),
            .I(N__47240));
    ClkMux I__11291 (
            .O(N__47683),
            .I(N__47240));
    ClkMux I__11290 (
            .O(N__47682),
            .I(N__47240));
    ClkMux I__11289 (
            .O(N__47681),
            .I(N__47240));
    ClkMux I__11288 (
            .O(N__47680),
            .I(N__47240));
    ClkMux I__11287 (
            .O(N__47679),
            .I(N__47240));
    ClkMux I__11286 (
            .O(N__47678),
            .I(N__47240));
    ClkMux I__11285 (
            .O(N__47677),
            .I(N__47240));
    ClkMux I__11284 (
            .O(N__47676),
            .I(N__47240));
    ClkMux I__11283 (
            .O(N__47675),
            .I(N__47240));
    ClkMux I__11282 (
            .O(N__47674),
            .I(N__47240));
    ClkMux I__11281 (
            .O(N__47673),
            .I(N__47240));
    ClkMux I__11280 (
            .O(N__47672),
            .I(N__47240));
    ClkMux I__11279 (
            .O(N__47671),
            .I(N__47240));
    ClkMux I__11278 (
            .O(N__47670),
            .I(N__47240));
    ClkMux I__11277 (
            .O(N__47669),
            .I(N__47240));
    ClkMux I__11276 (
            .O(N__47668),
            .I(N__47240));
    ClkMux I__11275 (
            .O(N__47667),
            .I(N__47240));
    ClkMux I__11274 (
            .O(N__47666),
            .I(N__47240));
    ClkMux I__11273 (
            .O(N__47665),
            .I(N__47240));
    ClkMux I__11272 (
            .O(N__47664),
            .I(N__47240));
    ClkMux I__11271 (
            .O(N__47663),
            .I(N__47240));
    ClkMux I__11270 (
            .O(N__47662),
            .I(N__47240));
    ClkMux I__11269 (
            .O(N__47661),
            .I(N__47240));
    ClkMux I__11268 (
            .O(N__47660),
            .I(N__47240));
    ClkMux I__11267 (
            .O(N__47659),
            .I(N__47240));
    ClkMux I__11266 (
            .O(N__47658),
            .I(N__47240));
    ClkMux I__11265 (
            .O(N__47657),
            .I(N__47240));
    ClkMux I__11264 (
            .O(N__47656),
            .I(N__47240));
    ClkMux I__11263 (
            .O(N__47655),
            .I(N__47240));
    ClkMux I__11262 (
            .O(N__47654),
            .I(N__47240));
    ClkMux I__11261 (
            .O(N__47653),
            .I(N__47240));
    ClkMux I__11260 (
            .O(N__47652),
            .I(N__47240));
    ClkMux I__11259 (
            .O(N__47651),
            .I(N__47240));
    ClkMux I__11258 (
            .O(N__47650),
            .I(N__47240));
    ClkMux I__11257 (
            .O(N__47649),
            .I(N__47240));
    ClkMux I__11256 (
            .O(N__47648),
            .I(N__47240));
    ClkMux I__11255 (
            .O(N__47647),
            .I(N__47240));
    ClkMux I__11254 (
            .O(N__47646),
            .I(N__47240));
    ClkMux I__11253 (
            .O(N__47645),
            .I(N__47240));
    ClkMux I__11252 (
            .O(N__47644),
            .I(N__47240));
    ClkMux I__11251 (
            .O(N__47643),
            .I(N__47240));
    ClkMux I__11250 (
            .O(N__47642),
            .I(N__47240));
    ClkMux I__11249 (
            .O(N__47641),
            .I(N__47240));
    ClkMux I__11248 (
            .O(N__47640),
            .I(N__47240));
    ClkMux I__11247 (
            .O(N__47639),
            .I(N__47240));
    ClkMux I__11246 (
            .O(N__47638),
            .I(N__47240));
    ClkMux I__11245 (
            .O(N__47637),
            .I(N__47240));
    ClkMux I__11244 (
            .O(N__47636),
            .I(N__47240));
    ClkMux I__11243 (
            .O(N__47635),
            .I(N__47240));
    ClkMux I__11242 (
            .O(N__47634),
            .I(N__47240));
    ClkMux I__11241 (
            .O(N__47633),
            .I(N__47240));
    ClkMux I__11240 (
            .O(N__47632),
            .I(N__47240));
    ClkMux I__11239 (
            .O(N__47631),
            .I(N__47240));
    ClkMux I__11238 (
            .O(N__47630),
            .I(N__47240));
    ClkMux I__11237 (
            .O(N__47629),
            .I(N__47240));
    ClkMux I__11236 (
            .O(N__47628),
            .I(N__47240));
    ClkMux I__11235 (
            .O(N__47627),
            .I(N__47240));
    ClkMux I__11234 (
            .O(N__47626),
            .I(N__47240));
    ClkMux I__11233 (
            .O(N__47625),
            .I(N__47240));
    ClkMux I__11232 (
            .O(N__47624),
            .I(N__47240));
    ClkMux I__11231 (
            .O(N__47623),
            .I(N__47240));
    ClkMux I__11230 (
            .O(N__47622),
            .I(N__47240));
    ClkMux I__11229 (
            .O(N__47621),
            .I(N__47240));
    ClkMux I__11228 (
            .O(N__47620),
            .I(N__47240));
    ClkMux I__11227 (
            .O(N__47619),
            .I(N__47240));
    ClkMux I__11226 (
            .O(N__47618),
            .I(N__47240));
    ClkMux I__11225 (
            .O(N__47617),
            .I(N__47240));
    ClkMux I__11224 (
            .O(N__47616),
            .I(N__47240));
    ClkMux I__11223 (
            .O(N__47615),
            .I(N__47240));
    ClkMux I__11222 (
            .O(N__47614),
            .I(N__47240));
    ClkMux I__11221 (
            .O(N__47613),
            .I(N__47240));
    ClkMux I__11220 (
            .O(N__47612),
            .I(N__47240));
    ClkMux I__11219 (
            .O(N__47611),
            .I(N__47240));
    ClkMux I__11218 (
            .O(N__47610),
            .I(N__47240));
    ClkMux I__11217 (
            .O(N__47609),
            .I(N__47240));
    ClkMux I__11216 (
            .O(N__47608),
            .I(N__47240));
    ClkMux I__11215 (
            .O(N__47607),
            .I(N__47240));
    ClkMux I__11214 (
            .O(N__47606),
            .I(N__47240));
    ClkMux I__11213 (
            .O(N__47605),
            .I(N__47240));
    ClkMux I__11212 (
            .O(N__47604),
            .I(N__47240));
    ClkMux I__11211 (
            .O(N__47603),
            .I(N__47240));
    ClkMux I__11210 (
            .O(N__47602),
            .I(N__47240));
    ClkMux I__11209 (
            .O(N__47601),
            .I(N__47240));
    ClkMux I__11208 (
            .O(N__47600),
            .I(N__47240));
    ClkMux I__11207 (
            .O(N__47599),
            .I(N__47240));
    ClkMux I__11206 (
            .O(N__47598),
            .I(N__47240));
    ClkMux I__11205 (
            .O(N__47597),
            .I(N__47240));
    ClkMux I__11204 (
            .O(N__47596),
            .I(N__47240));
    ClkMux I__11203 (
            .O(N__47595),
            .I(N__47240));
    ClkMux I__11202 (
            .O(N__47594),
            .I(N__47240));
    ClkMux I__11201 (
            .O(N__47593),
            .I(N__47240));
    ClkMux I__11200 (
            .O(N__47592),
            .I(N__47240));
    ClkMux I__11199 (
            .O(N__47591),
            .I(N__47240));
    ClkMux I__11198 (
            .O(N__47590),
            .I(N__47240));
    ClkMux I__11197 (
            .O(N__47589),
            .I(N__47240));
    ClkMux I__11196 (
            .O(N__47588),
            .I(N__47240));
    ClkMux I__11195 (
            .O(N__47587),
            .I(N__47240));
    ClkMux I__11194 (
            .O(N__47586),
            .I(N__47240));
    ClkMux I__11193 (
            .O(N__47585),
            .I(N__47240));
    ClkMux I__11192 (
            .O(N__47584),
            .I(N__47240));
    ClkMux I__11191 (
            .O(N__47583),
            .I(N__47240));
    ClkMux I__11190 (
            .O(N__47582),
            .I(N__47240));
    ClkMux I__11189 (
            .O(N__47581),
            .I(N__47240));
    ClkMux I__11188 (
            .O(N__47580),
            .I(N__47240));
    ClkMux I__11187 (
            .O(N__47579),
            .I(N__47240));
    ClkMux I__11186 (
            .O(N__47578),
            .I(N__47240));
    ClkMux I__11185 (
            .O(N__47577),
            .I(N__47240));
    ClkMux I__11184 (
            .O(N__47576),
            .I(N__47240));
    ClkMux I__11183 (
            .O(N__47575),
            .I(N__47240));
    ClkMux I__11182 (
            .O(N__47574),
            .I(N__47240));
    ClkMux I__11181 (
            .O(N__47573),
            .I(N__47240));
    ClkMux I__11180 (
            .O(N__47572),
            .I(N__47240));
    ClkMux I__11179 (
            .O(N__47571),
            .I(N__47240));
    ClkMux I__11178 (
            .O(N__47570),
            .I(N__47240));
    ClkMux I__11177 (
            .O(N__47569),
            .I(N__47240));
    ClkMux I__11176 (
            .O(N__47568),
            .I(N__47240));
    ClkMux I__11175 (
            .O(N__47567),
            .I(N__47240));
    ClkMux I__11174 (
            .O(N__47566),
            .I(N__47240));
    ClkMux I__11173 (
            .O(N__47565),
            .I(N__47240));
    ClkMux I__11172 (
            .O(N__47564),
            .I(N__47240));
    ClkMux I__11171 (
            .O(N__47563),
            .I(N__47240));
    ClkMux I__11170 (
            .O(N__47562),
            .I(N__47240));
    ClkMux I__11169 (
            .O(N__47561),
            .I(N__47240));
    ClkMux I__11168 (
            .O(N__47560),
            .I(N__47240));
    ClkMux I__11167 (
            .O(N__47559),
            .I(N__47240));
    ClkMux I__11166 (
            .O(N__47558),
            .I(N__47240));
    ClkMux I__11165 (
            .O(N__47557),
            .I(N__47240));
    ClkMux I__11164 (
            .O(N__47556),
            .I(N__47240));
    ClkMux I__11163 (
            .O(N__47555),
            .I(N__47240));
    ClkMux I__11162 (
            .O(N__47554),
            .I(N__47240));
    ClkMux I__11161 (
            .O(N__47553),
            .I(N__47240));
    ClkMux I__11160 (
            .O(N__47552),
            .I(N__47240));
    ClkMux I__11159 (
            .O(N__47551),
            .I(N__47240));
    ClkMux I__11158 (
            .O(N__47550),
            .I(N__47240));
    ClkMux I__11157 (
            .O(N__47549),
            .I(N__47240));
    GlobalMux I__11156 (
            .O(N__47240),
            .I(clk_100mhz_0));
    CEMux I__11155 (
            .O(N__47237),
            .I(N__47233));
    CEMux I__11154 (
            .O(N__47236),
            .I(N__47230));
    LocalMux I__11153 (
            .O(N__47233),
            .I(N__47224));
    LocalMux I__11152 (
            .O(N__47230),
            .I(N__47224));
    CEMux I__11151 (
            .O(N__47229),
            .I(N__47221));
    Span4Mux_v I__11150 (
            .O(N__47224),
            .I(N__47216));
    LocalMux I__11149 (
            .O(N__47221),
            .I(N__47213));
    CEMux I__11148 (
            .O(N__47220),
            .I(N__47210));
    CEMux I__11147 (
            .O(N__47219),
            .I(N__47205));
    Span4Mux_h I__11146 (
            .O(N__47216),
            .I(N__47195));
    Span4Mux_v I__11145 (
            .O(N__47213),
            .I(N__47195));
    LocalMux I__11144 (
            .O(N__47210),
            .I(N__47195));
    CEMux I__11143 (
            .O(N__47209),
            .I(N__47192));
    CEMux I__11142 (
            .O(N__47208),
            .I(N__47185));
    LocalMux I__11141 (
            .O(N__47205),
            .I(N__47182));
    CEMux I__11140 (
            .O(N__47204),
            .I(N__47179));
    CEMux I__11139 (
            .O(N__47203),
            .I(N__47176));
    CEMux I__11138 (
            .O(N__47202),
            .I(N__47173));
    Span4Mux_v I__11137 (
            .O(N__47195),
            .I(N__47166));
    LocalMux I__11136 (
            .O(N__47192),
            .I(N__47166));
    InMux I__11135 (
            .O(N__47191),
            .I(N__47147));
    InMux I__11134 (
            .O(N__47190),
            .I(N__47140));
    InMux I__11133 (
            .O(N__47189),
            .I(N__47140));
    InMux I__11132 (
            .O(N__47188),
            .I(N__47140));
    LocalMux I__11131 (
            .O(N__47185),
            .I(N__47137));
    Span4Mux_h I__11130 (
            .O(N__47182),
            .I(N__47134));
    LocalMux I__11129 (
            .O(N__47179),
            .I(N__47131));
    LocalMux I__11128 (
            .O(N__47176),
            .I(N__47126));
    LocalMux I__11127 (
            .O(N__47173),
            .I(N__47126));
    CEMux I__11126 (
            .O(N__47172),
            .I(N__47123));
    CEMux I__11125 (
            .O(N__47171),
            .I(N__47120));
    Span4Mux_v I__11124 (
            .O(N__47166),
            .I(N__47110));
    InMux I__11123 (
            .O(N__47165),
            .I(N__47101));
    InMux I__11122 (
            .O(N__47164),
            .I(N__47101));
    InMux I__11121 (
            .O(N__47163),
            .I(N__47101));
    InMux I__11120 (
            .O(N__47162),
            .I(N__47101));
    InMux I__11119 (
            .O(N__47161),
            .I(N__47092));
    InMux I__11118 (
            .O(N__47160),
            .I(N__47092));
    InMux I__11117 (
            .O(N__47159),
            .I(N__47092));
    InMux I__11116 (
            .O(N__47158),
            .I(N__47092));
    InMux I__11115 (
            .O(N__47157),
            .I(N__47083));
    InMux I__11114 (
            .O(N__47156),
            .I(N__47083));
    InMux I__11113 (
            .O(N__47155),
            .I(N__47083));
    InMux I__11112 (
            .O(N__47154),
            .I(N__47083));
    InMux I__11111 (
            .O(N__47153),
            .I(N__47074));
    InMux I__11110 (
            .O(N__47152),
            .I(N__47074));
    InMux I__11109 (
            .O(N__47151),
            .I(N__47074));
    InMux I__11108 (
            .O(N__47150),
            .I(N__47074));
    LocalMux I__11107 (
            .O(N__47147),
            .I(N__47071));
    LocalMux I__11106 (
            .O(N__47140),
            .I(N__47062));
    Span4Mux_v I__11105 (
            .O(N__47137),
            .I(N__47062));
    Span4Mux_v I__11104 (
            .O(N__47134),
            .I(N__47053));
    Span4Mux_v I__11103 (
            .O(N__47131),
            .I(N__47053));
    Span4Mux_h I__11102 (
            .O(N__47126),
            .I(N__47053));
    LocalMux I__11101 (
            .O(N__47123),
            .I(N__47053));
    LocalMux I__11100 (
            .O(N__47120),
            .I(N__47050));
    InMux I__11099 (
            .O(N__47119),
            .I(N__47043));
    InMux I__11098 (
            .O(N__47118),
            .I(N__47043));
    InMux I__11097 (
            .O(N__47117),
            .I(N__47043));
    InMux I__11096 (
            .O(N__47116),
            .I(N__47034));
    InMux I__11095 (
            .O(N__47115),
            .I(N__47034));
    InMux I__11094 (
            .O(N__47114),
            .I(N__47034));
    InMux I__11093 (
            .O(N__47113),
            .I(N__47034));
    Span4Mux_v I__11092 (
            .O(N__47110),
            .I(N__47029));
    LocalMux I__11091 (
            .O(N__47101),
            .I(N__47029));
    LocalMux I__11090 (
            .O(N__47092),
            .I(N__47026));
    LocalMux I__11089 (
            .O(N__47083),
            .I(N__47019));
    LocalMux I__11088 (
            .O(N__47074),
            .I(N__47019));
    Span4Mux_h I__11087 (
            .O(N__47071),
            .I(N__47019));
    InMux I__11086 (
            .O(N__47070),
            .I(N__47010));
    InMux I__11085 (
            .O(N__47069),
            .I(N__47010));
    InMux I__11084 (
            .O(N__47068),
            .I(N__47010));
    InMux I__11083 (
            .O(N__47067),
            .I(N__47010));
    Span4Mux_h I__11082 (
            .O(N__47062),
            .I(N__47005));
    Span4Mux_v I__11081 (
            .O(N__47053),
            .I(N__47005));
    Span4Mux_v I__11080 (
            .O(N__47050),
            .I(N__46998));
    LocalMux I__11079 (
            .O(N__47043),
            .I(N__46998));
    LocalMux I__11078 (
            .O(N__47034),
            .I(N__46998));
    Span4Mux_v I__11077 (
            .O(N__47029),
            .I(N__46993));
    Span4Mux_v I__11076 (
            .O(N__47026),
            .I(N__46993));
    Span4Mux_h I__11075 (
            .O(N__47019),
            .I(N__46990));
    LocalMux I__11074 (
            .O(N__47010),
            .I(N__46987));
    Span4Mux_h I__11073 (
            .O(N__47005),
            .I(N__46984));
    Span4Mux_h I__11072 (
            .O(N__46998),
            .I(N__46981));
    Span4Mux_h I__11071 (
            .O(N__46993),
            .I(N__46978));
    Span4Mux_h I__11070 (
            .O(N__46990),
            .I(N__46975));
    Span4Mux_h I__11069 (
            .O(N__46987),
            .I(N__46970));
    Span4Mux_s2_h I__11068 (
            .O(N__46984),
            .I(N__46970));
    Odrv4 I__11067 (
            .O(N__46981),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11066 (
            .O(N__46978),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11065 (
            .O(N__46975),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    Odrv4 I__11064 (
            .O(N__46970),
            .I(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ));
    InMux I__11063 (
            .O(N__46961),
            .I(N__46955));
    InMux I__11062 (
            .O(N__46960),
            .I(N__46950));
    InMux I__11061 (
            .O(N__46959),
            .I(N__46950));
    InMux I__11060 (
            .O(N__46958),
            .I(N__46947));
    LocalMux I__11059 (
            .O(N__46955),
            .I(N__46944));
    LocalMux I__11058 (
            .O(N__46950),
            .I(N__46941));
    LocalMux I__11057 (
            .O(N__46947),
            .I(N__46933));
    Glb2LocalMux I__11056 (
            .O(N__46944),
            .I(N__46466));
    Glb2LocalMux I__11055 (
            .O(N__46941),
            .I(N__46466));
    SRMux I__11054 (
            .O(N__46940),
            .I(N__46466));
    SRMux I__11053 (
            .O(N__46939),
            .I(N__46466));
    SRMux I__11052 (
            .O(N__46938),
            .I(N__46466));
    SRMux I__11051 (
            .O(N__46937),
            .I(N__46466));
    SRMux I__11050 (
            .O(N__46936),
            .I(N__46466));
    Glb2LocalMux I__11049 (
            .O(N__46933),
            .I(N__46466));
    SRMux I__11048 (
            .O(N__46932),
            .I(N__46466));
    SRMux I__11047 (
            .O(N__46931),
            .I(N__46466));
    SRMux I__11046 (
            .O(N__46930),
            .I(N__46466));
    SRMux I__11045 (
            .O(N__46929),
            .I(N__46466));
    SRMux I__11044 (
            .O(N__46928),
            .I(N__46466));
    SRMux I__11043 (
            .O(N__46927),
            .I(N__46466));
    SRMux I__11042 (
            .O(N__46926),
            .I(N__46466));
    SRMux I__11041 (
            .O(N__46925),
            .I(N__46466));
    SRMux I__11040 (
            .O(N__46924),
            .I(N__46466));
    SRMux I__11039 (
            .O(N__46923),
            .I(N__46466));
    SRMux I__11038 (
            .O(N__46922),
            .I(N__46466));
    SRMux I__11037 (
            .O(N__46921),
            .I(N__46466));
    SRMux I__11036 (
            .O(N__46920),
            .I(N__46466));
    SRMux I__11035 (
            .O(N__46919),
            .I(N__46466));
    SRMux I__11034 (
            .O(N__46918),
            .I(N__46466));
    SRMux I__11033 (
            .O(N__46917),
            .I(N__46466));
    SRMux I__11032 (
            .O(N__46916),
            .I(N__46466));
    SRMux I__11031 (
            .O(N__46915),
            .I(N__46466));
    SRMux I__11030 (
            .O(N__46914),
            .I(N__46466));
    SRMux I__11029 (
            .O(N__46913),
            .I(N__46466));
    SRMux I__11028 (
            .O(N__46912),
            .I(N__46466));
    SRMux I__11027 (
            .O(N__46911),
            .I(N__46466));
    SRMux I__11026 (
            .O(N__46910),
            .I(N__46466));
    SRMux I__11025 (
            .O(N__46909),
            .I(N__46466));
    SRMux I__11024 (
            .O(N__46908),
            .I(N__46466));
    SRMux I__11023 (
            .O(N__46907),
            .I(N__46466));
    SRMux I__11022 (
            .O(N__46906),
            .I(N__46466));
    SRMux I__11021 (
            .O(N__46905),
            .I(N__46466));
    SRMux I__11020 (
            .O(N__46904),
            .I(N__46466));
    SRMux I__11019 (
            .O(N__46903),
            .I(N__46466));
    SRMux I__11018 (
            .O(N__46902),
            .I(N__46466));
    SRMux I__11017 (
            .O(N__46901),
            .I(N__46466));
    SRMux I__11016 (
            .O(N__46900),
            .I(N__46466));
    SRMux I__11015 (
            .O(N__46899),
            .I(N__46466));
    SRMux I__11014 (
            .O(N__46898),
            .I(N__46466));
    SRMux I__11013 (
            .O(N__46897),
            .I(N__46466));
    SRMux I__11012 (
            .O(N__46896),
            .I(N__46466));
    SRMux I__11011 (
            .O(N__46895),
            .I(N__46466));
    SRMux I__11010 (
            .O(N__46894),
            .I(N__46466));
    SRMux I__11009 (
            .O(N__46893),
            .I(N__46466));
    SRMux I__11008 (
            .O(N__46892),
            .I(N__46466));
    SRMux I__11007 (
            .O(N__46891),
            .I(N__46466));
    SRMux I__11006 (
            .O(N__46890),
            .I(N__46466));
    SRMux I__11005 (
            .O(N__46889),
            .I(N__46466));
    SRMux I__11004 (
            .O(N__46888),
            .I(N__46466));
    SRMux I__11003 (
            .O(N__46887),
            .I(N__46466));
    SRMux I__11002 (
            .O(N__46886),
            .I(N__46466));
    SRMux I__11001 (
            .O(N__46885),
            .I(N__46466));
    SRMux I__11000 (
            .O(N__46884),
            .I(N__46466));
    SRMux I__10999 (
            .O(N__46883),
            .I(N__46466));
    SRMux I__10998 (
            .O(N__46882),
            .I(N__46466));
    SRMux I__10997 (
            .O(N__46881),
            .I(N__46466));
    SRMux I__10996 (
            .O(N__46880),
            .I(N__46466));
    SRMux I__10995 (
            .O(N__46879),
            .I(N__46466));
    SRMux I__10994 (
            .O(N__46878),
            .I(N__46466));
    SRMux I__10993 (
            .O(N__46877),
            .I(N__46466));
    SRMux I__10992 (
            .O(N__46876),
            .I(N__46466));
    SRMux I__10991 (
            .O(N__46875),
            .I(N__46466));
    SRMux I__10990 (
            .O(N__46874),
            .I(N__46466));
    SRMux I__10989 (
            .O(N__46873),
            .I(N__46466));
    SRMux I__10988 (
            .O(N__46872),
            .I(N__46466));
    SRMux I__10987 (
            .O(N__46871),
            .I(N__46466));
    SRMux I__10986 (
            .O(N__46870),
            .I(N__46466));
    SRMux I__10985 (
            .O(N__46869),
            .I(N__46466));
    SRMux I__10984 (
            .O(N__46868),
            .I(N__46466));
    SRMux I__10983 (
            .O(N__46867),
            .I(N__46466));
    SRMux I__10982 (
            .O(N__46866),
            .I(N__46466));
    SRMux I__10981 (
            .O(N__46865),
            .I(N__46466));
    SRMux I__10980 (
            .O(N__46864),
            .I(N__46466));
    SRMux I__10979 (
            .O(N__46863),
            .I(N__46466));
    SRMux I__10978 (
            .O(N__46862),
            .I(N__46466));
    SRMux I__10977 (
            .O(N__46861),
            .I(N__46466));
    SRMux I__10976 (
            .O(N__46860),
            .I(N__46466));
    SRMux I__10975 (
            .O(N__46859),
            .I(N__46466));
    SRMux I__10974 (
            .O(N__46858),
            .I(N__46466));
    SRMux I__10973 (
            .O(N__46857),
            .I(N__46466));
    SRMux I__10972 (
            .O(N__46856),
            .I(N__46466));
    SRMux I__10971 (
            .O(N__46855),
            .I(N__46466));
    SRMux I__10970 (
            .O(N__46854),
            .I(N__46466));
    SRMux I__10969 (
            .O(N__46853),
            .I(N__46466));
    SRMux I__10968 (
            .O(N__46852),
            .I(N__46466));
    SRMux I__10967 (
            .O(N__46851),
            .I(N__46466));
    SRMux I__10966 (
            .O(N__46850),
            .I(N__46466));
    SRMux I__10965 (
            .O(N__46849),
            .I(N__46466));
    SRMux I__10964 (
            .O(N__46848),
            .I(N__46466));
    SRMux I__10963 (
            .O(N__46847),
            .I(N__46466));
    SRMux I__10962 (
            .O(N__46846),
            .I(N__46466));
    SRMux I__10961 (
            .O(N__46845),
            .I(N__46466));
    SRMux I__10960 (
            .O(N__46844),
            .I(N__46466));
    SRMux I__10959 (
            .O(N__46843),
            .I(N__46466));
    SRMux I__10958 (
            .O(N__46842),
            .I(N__46466));
    SRMux I__10957 (
            .O(N__46841),
            .I(N__46466));
    SRMux I__10956 (
            .O(N__46840),
            .I(N__46466));
    SRMux I__10955 (
            .O(N__46839),
            .I(N__46466));
    SRMux I__10954 (
            .O(N__46838),
            .I(N__46466));
    SRMux I__10953 (
            .O(N__46837),
            .I(N__46466));
    SRMux I__10952 (
            .O(N__46836),
            .I(N__46466));
    SRMux I__10951 (
            .O(N__46835),
            .I(N__46466));
    SRMux I__10950 (
            .O(N__46834),
            .I(N__46466));
    SRMux I__10949 (
            .O(N__46833),
            .I(N__46466));
    SRMux I__10948 (
            .O(N__46832),
            .I(N__46466));
    SRMux I__10947 (
            .O(N__46831),
            .I(N__46466));
    SRMux I__10946 (
            .O(N__46830),
            .I(N__46466));
    SRMux I__10945 (
            .O(N__46829),
            .I(N__46466));
    SRMux I__10944 (
            .O(N__46828),
            .I(N__46466));
    SRMux I__10943 (
            .O(N__46827),
            .I(N__46466));
    SRMux I__10942 (
            .O(N__46826),
            .I(N__46466));
    SRMux I__10941 (
            .O(N__46825),
            .I(N__46466));
    SRMux I__10940 (
            .O(N__46824),
            .I(N__46466));
    SRMux I__10939 (
            .O(N__46823),
            .I(N__46466));
    SRMux I__10938 (
            .O(N__46822),
            .I(N__46466));
    SRMux I__10937 (
            .O(N__46821),
            .I(N__46466));
    SRMux I__10936 (
            .O(N__46820),
            .I(N__46466));
    SRMux I__10935 (
            .O(N__46819),
            .I(N__46466));
    SRMux I__10934 (
            .O(N__46818),
            .I(N__46466));
    SRMux I__10933 (
            .O(N__46817),
            .I(N__46466));
    SRMux I__10932 (
            .O(N__46816),
            .I(N__46466));
    SRMux I__10931 (
            .O(N__46815),
            .I(N__46466));
    SRMux I__10930 (
            .O(N__46814),
            .I(N__46466));
    SRMux I__10929 (
            .O(N__46813),
            .I(N__46466));
    SRMux I__10928 (
            .O(N__46812),
            .I(N__46466));
    SRMux I__10927 (
            .O(N__46811),
            .I(N__46466));
    SRMux I__10926 (
            .O(N__46810),
            .I(N__46466));
    SRMux I__10925 (
            .O(N__46809),
            .I(N__46466));
    SRMux I__10924 (
            .O(N__46808),
            .I(N__46466));
    SRMux I__10923 (
            .O(N__46807),
            .I(N__46466));
    SRMux I__10922 (
            .O(N__46806),
            .I(N__46466));
    SRMux I__10921 (
            .O(N__46805),
            .I(N__46466));
    SRMux I__10920 (
            .O(N__46804),
            .I(N__46466));
    SRMux I__10919 (
            .O(N__46803),
            .I(N__46466));
    SRMux I__10918 (
            .O(N__46802),
            .I(N__46466));
    SRMux I__10917 (
            .O(N__46801),
            .I(N__46466));
    SRMux I__10916 (
            .O(N__46800),
            .I(N__46466));
    SRMux I__10915 (
            .O(N__46799),
            .I(N__46466));
    SRMux I__10914 (
            .O(N__46798),
            .I(N__46466));
    SRMux I__10913 (
            .O(N__46797),
            .I(N__46466));
    SRMux I__10912 (
            .O(N__46796),
            .I(N__46466));
    SRMux I__10911 (
            .O(N__46795),
            .I(N__46466));
    SRMux I__10910 (
            .O(N__46794),
            .I(N__46466));
    SRMux I__10909 (
            .O(N__46793),
            .I(N__46466));
    SRMux I__10908 (
            .O(N__46792),
            .I(N__46466));
    SRMux I__10907 (
            .O(N__46791),
            .I(N__46466));
    SRMux I__10906 (
            .O(N__46790),
            .I(N__46466));
    SRMux I__10905 (
            .O(N__46789),
            .I(N__46466));
    SRMux I__10904 (
            .O(N__46788),
            .I(N__46466));
    SRMux I__10903 (
            .O(N__46787),
            .I(N__46466));
    SRMux I__10902 (
            .O(N__46786),
            .I(N__46466));
    SRMux I__10901 (
            .O(N__46785),
            .I(N__46466));
    SRMux I__10900 (
            .O(N__46784),
            .I(N__46466));
    SRMux I__10899 (
            .O(N__46783),
            .I(N__46466));
    GlobalMux I__10898 (
            .O(N__46466),
            .I(N__46463));
    gio2CtrlBuf I__10897 (
            .O(N__46463),
            .I(red_c_g));
    CascadeMux I__10896 (
            .O(N__46460),
            .I(N__46457));
    InMux I__10895 (
            .O(N__46457),
            .I(N__46454));
    LocalMux I__10894 (
            .O(N__46454),
            .I(N__46451));
    Span4Mux_h I__10893 (
            .O(N__46451),
            .I(N__46448));
    Odrv4 I__10892 (
            .O(N__46448),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt24 ));
    InMux I__10891 (
            .O(N__46445),
            .I(N__46439));
    InMux I__10890 (
            .O(N__46444),
            .I(N__46439));
    LocalMux I__10889 (
            .O(N__46439),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    InMux I__10888 (
            .O(N__46436),
            .I(N__46429));
    InMux I__10887 (
            .O(N__46435),
            .I(N__46429));
    InMux I__10886 (
            .O(N__46434),
            .I(N__46426));
    LocalMux I__10885 (
            .O(N__46429),
            .I(N__46423));
    LocalMux I__10884 (
            .O(N__46426),
            .I(N__46418));
    Span4Mux_h I__10883 (
            .O(N__46423),
            .I(N__46418));
    Odrv4 I__10882 (
            .O(N__46418),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    CascadeMux I__10881 (
            .O(N__46415),
            .I(N__46411));
    CascadeMux I__10880 (
            .O(N__46414),
            .I(N__46408));
    InMux I__10879 (
            .O(N__46411),
            .I(N__46403));
    InMux I__10878 (
            .O(N__46408),
            .I(N__46403));
    LocalMux I__10877 (
            .O(N__46403),
            .I(N__46399));
    InMux I__10876 (
            .O(N__46402),
            .I(N__46396));
    Span4Mux_h I__10875 (
            .O(N__46399),
            .I(N__46393));
    LocalMux I__10874 (
            .O(N__46396),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__10873 (
            .O(N__46393),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__10872 (
            .O(N__46388),
            .I(N__46382));
    InMux I__10871 (
            .O(N__46387),
            .I(N__46382));
    LocalMux I__10870 (
            .O(N__46382),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ));
    InMux I__10869 (
            .O(N__46379),
            .I(N__46376));
    LocalMux I__10868 (
            .O(N__46376),
            .I(N__46373));
    Odrv12 I__10867 (
            .O(N__46373),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ));
    CascadeMux I__10866 (
            .O(N__46370),
            .I(N__46367));
    InMux I__10865 (
            .O(N__46367),
            .I(N__46362));
    InMux I__10864 (
            .O(N__46366),
            .I(N__46359));
    InMux I__10863 (
            .O(N__46365),
            .I(N__46356));
    LocalMux I__10862 (
            .O(N__46362),
            .I(N__46351));
    LocalMux I__10861 (
            .O(N__46359),
            .I(N__46351));
    LocalMux I__10860 (
            .O(N__46356),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv12 I__10859 (
            .O(N__46351),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__10858 (
            .O(N__46346),
            .I(N__46342));
    InMux I__10857 (
            .O(N__46345),
            .I(N__46339));
    LocalMux I__10856 (
            .O(N__46342),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    LocalMux I__10855 (
            .O(N__46339),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    CascadeMux I__10854 (
            .O(N__46334),
            .I(N__46331));
    InMux I__10853 (
            .O(N__46331),
            .I(N__46326));
    InMux I__10852 (
            .O(N__46330),
            .I(N__46323));
    InMux I__10851 (
            .O(N__46329),
            .I(N__46320));
    LocalMux I__10850 (
            .O(N__46326),
            .I(N__46317));
    LocalMux I__10849 (
            .O(N__46323),
            .I(N__46314));
    LocalMux I__10848 (
            .O(N__46320),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv12 I__10847 (
            .O(N__46317),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__10846 (
            .O(N__46314),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__10845 (
            .O(N__46307),
            .I(N__46303));
    InMux I__10844 (
            .O(N__46306),
            .I(N__46300));
    LocalMux I__10843 (
            .O(N__46303),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    LocalMux I__10842 (
            .O(N__46300),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    CascadeMux I__10841 (
            .O(N__46295),
            .I(N__46292));
    InMux I__10840 (
            .O(N__46292),
            .I(N__46289));
    LocalMux I__10839 (
            .O(N__46289),
            .I(N__46286));
    Odrv12 I__10838 (
            .O(N__46286),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ));
    InMux I__10837 (
            .O(N__46283),
            .I(N__46280));
    LocalMux I__10836 (
            .O(N__46280),
            .I(N__46277));
    Span4Mux_v I__10835 (
            .O(N__46277),
            .I(N__46274));
    Sp12to4 I__10834 (
            .O(N__46274),
            .I(N__46271));
    Span12Mux_h I__10833 (
            .O(N__46271),
            .I(N__46267));
    InMux I__10832 (
            .O(N__46270),
            .I(N__46264));
    Odrv12 I__10831 (
            .O(N__46267),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    LocalMux I__10830 (
            .O(N__46264),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    CascadeMux I__10829 (
            .O(N__46259),
            .I(N__46256));
    InMux I__10828 (
            .O(N__46256),
            .I(N__46250));
    CascadeMux I__10827 (
            .O(N__46255),
            .I(N__46244));
    CascadeMux I__10826 (
            .O(N__46254),
            .I(N__46239));
    CascadeMux I__10825 (
            .O(N__46253),
            .I(N__46236));
    LocalMux I__10824 (
            .O(N__46250),
            .I(N__46228));
    InMux I__10823 (
            .O(N__46249),
            .I(N__46219));
    InMux I__10822 (
            .O(N__46248),
            .I(N__46219));
    InMux I__10821 (
            .O(N__46247),
            .I(N__46219));
    InMux I__10820 (
            .O(N__46244),
            .I(N__46219));
    InMux I__10819 (
            .O(N__46243),
            .I(N__46210));
    InMux I__10818 (
            .O(N__46242),
            .I(N__46210));
    InMux I__10817 (
            .O(N__46239),
            .I(N__46210));
    InMux I__10816 (
            .O(N__46236),
            .I(N__46210));
    InMux I__10815 (
            .O(N__46235),
            .I(N__46203));
    InMux I__10814 (
            .O(N__46234),
            .I(N__46203));
    InMux I__10813 (
            .O(N__46233),
            .I(N__46196));
    InMux I__10812 (
            .O(N__46232),
            .I(N__46196));
    InMux I__10811 (
            .O(N__46231),
            .I(N__46196));
    Span4Mux_v I__10810 (
            .O(N__46228),
            .I(N__46191));
    LocalMux I__10809 (
            .O(N__46219),
            .I(N__46191));
    LocalMux I__10808 (
            .O(N__46210),
            .I(N__46188));
    InMux I__10807 (
            .O(N__46209),
            .I(N__46185));
    CascadeMux I__10806 (
            .O(N__46208),
            .I(N__46166));
    LocalMux I__10805 (
            .O(N__46203),
            .I(N__46163));
    LocalMux I__10804 (
            .O(N__46196),
            .I(N__46160));
    Span4Mux_h I__10803 (
            .O(N__46191),
            .I(N__46155));
    Span4Mux_v I__10802 (
            .O(N__46188),
            .I(N__46155));
    LocalMux I__10801 (
            .O(N__46185),
            .I(N__46152));
    InMux I__10800 (
            .O(N__46184),
            .I(N__46135));
    InMux I__10799 (
            .O(N__46183),
            .I(N__46135));
    InMux I__10798 (
            .O(N__46182),
            .I(N__46135));
    InMux I__10797 (
            .O(N__46181),
            .I(N__46135));
    InMux I__10796 (
            .O(N__46180),
            .I(N__46135));
    InMux I__10795 (
            .O(N__46179),
            .I(N__46135));
    InMux I__10794 (
            .O(N__46178),
            .I(N__46135));
    InMux I__10793 (
            .O(N__46177),
            .I(N__46135));
    InMux I__10792 (
            .O(N__46176),
            .I(N__46120));
    InMux I__10791 (
            .O(N__46175),
            .I(N__46120));
    InMux I__10790 (
            .O(N__46174),
            .I(N__46120));
    InMux I__10789 (
            .O(N__46173),
            .I(N__46120));
    InMux I__10788 (
            .O(N__46172),
            .I(N__46120));
    InMux I__10787 (
            .O(N__46171),
            .I(N__46120));
    InMux I__10786 (
            .O(N__46170),
            .I(N__46120));
    InMux I__10785 (
            .O(N__46169),
            .I(N__46117));
    InMux I__10784 (
            .O(N__46166),
            .I(N__46114));
    Span4Mux_v I__10783 (
            .O(N__46163),
            .I(N__46111));
    Sp12to4 I__10782 (
            .O(N__46160),
            .I(N__46108));
    Span4Mux_h I__10781 (
            .O(N__46155),
            .I(N__46105));
    Sp12to4 I__10780 (
            .O(N__46152),
            .I(N__46098));
    LocalMux I__10779 (
            .O(N__46135),
            .I(N__46098));
    LocalMux I__10778 (
            .O(N__46120),
            .I(N__46098));
    LocalMux I__10777 (
            .O(N__46117),
            .I(N__46089));
    LocalMux I__10776 (
            .O(N__46114),
            .I(N__46089));
    Sp12to4 I__10775 (
            .O(N__46111),
            .I(N__46089));
    Span12Mux_s7_v I__10774 (
            .O(N__46108),
            .I(N__46089));
    Sp12to4 I__10773 (
            .O(N__46105),
            .I(N__46082));
    Span12Mux_s7_v I__10772 (
            .O(N__46098),
            .I(N__46082));
    Span12Mux_h I__10771 (
            .O(N__46089),
            .I(N__46082));
    Odrv12 I__10770 (
            .O(N__46082),
            .I(N_19_1));
    InMux I__10769 (
            .O(N__46079),
            .I(N__46076));
    LocalMux I__10768 (
            .O(N__46076),
            .I(N__46068));
    InMux I__10767 (
            .O(N__46075),
            .I(N__46065));
    CascadeMux I__10766 (
            .O(N__46074),
            .I(N__46061));
    CascadeMux I__10765 (
            .O(N__46073),
            .I(N__46058));
    CascadeMux I__10764 (
            .O(N__46072),
            .I(N__46054));
    CascadeMux I__10763 (
            .O(N__46071),
            .I(N__46051));
    Span12Mux_s7_v I__10762 (
            .O(N__46068),
            .I(N__46048));
    LocalMux I__10761 (
            .O(N__46065),
            .I(N__46045));
    InMux I__10760 (
            .O(N__46064),
            .I(N__46038));
    InMux I__10759 (
            .O(N__46061),
            .I(N__46038));
    InMux I__10758 (
            .O(N__46058),
            .I(N__46038));
    InMux I__10757 (
            .O(N__46057),
            .I(N__46031));
    InMux I__10756 (
            .O(N__46054),
            .I(N__46031));
    InMux I__10755 (
            .O(N__46051),
            .I(N__46031));
    Span12Mux_h I__10754 (
            .O(N__46048),
            .I(N__46028));
    Span4Mux_v I__10753 (
            .O(N__46045),
            .I(N__46021));
    LocalMux I__10752 (
            .O(N__46038),
            .I(N__46021));
    LocalMux I__10751 (
            .O(N__46031),
            .I(N__46021));
    Span12Mux_h I__10750 (
            .O(N__46028),
            .I(N__46018));
    Span4Mux_h I__10749 (
            .O(N__46021),
            .I(N__46015));
    Odrv12 I__10748 (
            .O(N__46018),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    Odrv4 I__10747 (
            .O(N__46015),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    CascadeMux I__10746 (
            .O(N__46010),
            .I(N__46007));
    InMux I__10745 (
            .O(N__46007),
            .I(N__46004));
    LocalMux I__10744 (
            .O(N__46004),
            .I(N__46001));
    Span12Mux_s7_h I__10743 (
            .O(N__46001),
            .I(N__45998));
    Span12Mux_h I__10742 (
            .O(N__45998),
            .I(N__45995));
    Odrv12 I__10741 (
            .O(N__45995),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    InMux I__10740 (
            .O(N__45992),
            .I(N__45986));
    InMux I__10739 (
            .O(N__45991),
            .I(N__45986));
    LocalMux I__10738 (
            .O(N__45986),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    CascadeMux I__10737 (
            .O(N__45983),
            .I(N__45980));
    InMux I__10736 (
            .O(N__45980),
            .I(N__45974));
    InMux I__10735 (
            .O(N__45979),
            .I(N__45974));
    LocalMux I__10734 (
            .O(N__45974),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    InMux I__10733 (
            .O(N__45971),
            .I(N__45967));
    InMux I__10732 (
            .O(N__45970),
            .I(N__45964));
    LocalMux I__10731 (
            .O(N__45967),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    LocalMux I__10730 (
            .O(N__45964),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    CEMux I__10729 (
            .O(N__45959),
            .I(N__45935));
    CEMux I__10728 (
            .O(N__45958),
            .I(N__45935));
    CEMux I__10727 (
            .O(N__45957),
            .I(N__45935));
    CEMux I__10726 (
            .O(N__45956),
            .I(N__45935));
    CEMux I__10725 (
            .O(N__45955),
            .I(N__45935));
    CEMux I__10724 (
            .O(N__45954),
            .I(N__45935));
    CEMux I__10723 (
            .O(N__45953),
            .I(N__45935));
    CEMux I__10722 (
            .O(N__45952),
            .I(N__45935));
    GlobalMux I__10721 (
            .O(N__45935),
            .I(N__45932));
    gio2CtrlBuf I__10720 (
            .O(N__45932),
            .I(\phase_controller_inst2.stoper_tr.un1_start_g ));
    InMux I__10719 (
            .O(N__45929),
            .I(N__45923));
    InMux I__10718 (
            .O(N__45928),
            .I(N__45920));
    InMux I__10717 (
            .O(N__45927),
            .I(N__45917));
    InMux I__10716 (
            .O(N__45926),
            .I(N__45914));
    LocalMux I__10715 (
            .O(N__45923),
            .I(N__45911));
    LocalMux I__10714 (
            .O(N__45920),
            .I(N__45906));
    LocalMux I__10713 (
            .O(N__45917),
            .I(N__45906));
    LocalMux I__10712 (
            .O(N__45914),
            .I(N__45903));
    Span4Mux_h I__10711 (
            .O(N__45911),
            .I(N__45900));
    Span4Mux_h I__10710 (
            .O(N__45906),
            .I(N__45895));
    Span4Mux_v I__10709 (
            .O(N__45903),
            .I(N__45895));
    Span4Mux_h I__10708 (
            .O(N__45900),
            .I(N__45892));
    Span4Mux_h I__10707 (
            .O(N__45895),
            .I(N__45889));
    Odrv4 I__10706 (
            .O(N__45892),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__10705 (
            .O(N__45889),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__10704 (
            .O(N__45884),
            .I(N__45879));
    InMux I__10703 (
            .O(N__45883),
            .I(N__45876));
    InMux I__10702 (
            .O(N__45882),
            .I(N__45873));
    LocalMux I__10701 (
            .O(N__45879),
            .I(N__45868));
    LocalMux I__10700 (
            .O(N__45876),
            .I(N__45868));
    LocalMux I__10699 (
            .O(N__45873),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv4 I__10698 (
            .O(N__45868),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    InMux I__10697 (
            .O(N__45863),
            .I(N__45859));
    InMux I__10696 (
            .O(N__45862),
            .I(N__45855));
    LocalMux I__10695 (
            .O(N__45859),
            .I(N__45852));
    InMux I__10694 (
            .O(N__45858),
            .I(N__45849));
    LocalMux I__10693 (
            .O(N__45855),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    Odrv4 I__10692 (
            .O(N__45852),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    LocalMux I__10691 (
            .O(N__45849),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__10690 (
            .O(N__45842),
            .I(N__45837));
    InMux I__10689 (
            .O(N__45841),
            .I(N__45834));
    CascadeMux I__10688 (
            .O(N__45840),
            .I(N__45831));
    LocalMux I__10687 (
            .O(N__45837),
            .I(N__45827));
    LocalMux I__10686 (
            .O(N__45834),
            .I(N__45824));
    InMux I__10685 (
            .O(N__45831),
            .I(N__45821));
    InMux I__10684 (
            .O(N__45830),
            .I(N__45818));
    Span4Mux_v I__10683 (
            .O(N__45827),
            .I(N__45815));
    Span4Mux_h I__10682 (
            .O(N__45824),
            .I(N__45812));
    LocalMux I__10681 (
            .O(N__45821),
            .I(N__45809));
    LocalMux I__10680 (
            .O(N__45818),
            .I(N__45806));
    Span4Mux_h I__10679 (
            .O(N__45815),
            .I(N__45803));
    Span4Mux_h I__10678 (
            .O(N__45812),
            .I(N__45800));
    Span12Mux_s11_v I__10677 (
            .O(N__45809),
            .I(N__45797));
    Odrv12 I__10676 (
            .O(N__45806),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv4 I__10675 (
            .O(N__45803),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv4 I__10674 (
            .O(N__45800),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv12 I__10673 (
            .O(N__45797),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__10672 (
            .O(N__45788),
            .I(N__45783));
    InMux I__10671 (
            .O(N__45787),
            .I(N__45780));
    InMux I__10670 (
            .O(N__45786),
            .I(N__45777));
    LocalMux I__10669 (
            .O(N__45783),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    LocalMux I__10668 (
            .O(N__45780),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    LocalMux I__10667 (
            .O(N__45777),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    InMux I__10666 (
            .O(N__45770),
            .I(N__45766));
    InMux I__10665 (
            .O(N__45769),
            .I(N__45763));
    LocalMux I__10664 (
            .O(N__45766),
            .I(N__45758));
    LocalMux I__10663 (
            .O(N__45763),
            .I(N__45758));
    Span4Mux_v I__10662 (
            .O(N__45758),
            .I(N__45753));
    InMux I__10661 (
            .O(N__45757),
            .I(N__45750));
    InMux I__10660 (
            .O(N__45756),
            .I(N__45747));
    Sp12to4 I__10659 (
            .O(N__45753),
            .I(N__45742));
    LocalMux I__10658 (
            .O(N__45750),
            .I(N__45742));
    LocalMux I__10657 (
            .O(N__45747),
            .I(N__45739));
    Span12Mux_s10_h I__10656 (
            .O(N__45742),
            .I(N__45736));
    Odrv12 I__10655 (
            .O(N__45739),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv12 I__10654 (
            .O(N__45736),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    CascadeMux I__10653 (
            .O(N__45731),
            .I(N__45728));
    InMux I__10652 (
            .O(N__45728),
            .I(N__45725));
    LocalMux I__10651 (
            .O(N__45725),
            .I(N__45722));
    Span4Mux_h I__10650 (
            .O(N__45722),
            .I(N__45719));
    Span4Mux_h I__10649 (
            .O(N__45719),
            .I(N__45716));
    Odrv4 I__10648 (
            .O(N__45716),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ));
    InMux I__10647 (
            .O(N__45713),
            .I(N__45709));
    InMux I__10646 (
            .O(N__45712),
            .I(N__45706));
    LocalMux I__10645 (
            .O(N__45709),
            .I(N__45699));
    LocalMux I__10644 (
            .O(N__45706),
            .I(N__45699));
    InMux I__10643 (
            .O(N__45705),
            .I(N__45696));
    InMux I__10642 (
            .O(N__45704),
            .I(N__45693));
    Span4Mux_v I__10641 (
            .O(N__45699),
            .I(N__45688));
    LocalMux I__10640 (
            .O(N__45696),
            .I(N__45688));
    LocalMux I__10639 (
            .O(N__45693),
            .I(N__45685));
    Span4Mux_h I__10638 (
            .O(N__45688),
            .I(N__45682));
    Span4Mux_h I__10637 (
            .O(N__45685),
            .I(N__45679));
    Span4Mux_v I__10636 (
            .O(N__45682),
            .I(N__45676));
    Span4Mux_v I__10635 (
            .O(N__45679),
            .I(N__45673));
    Odrv4 I__10634 (
            .O(N__45676),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__10633 (
            .O(N__45673),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__10632 (
            .O(N__45668),
            .I(N__45664));
    InMux I__10631 (
            .O(N__45667),
            .I(N__45660));
    LocalMux I__10630 (
            .O(N__45664),
            .I(N__45657));
    InMux I__10629 (
            .O(N__45663),
            .I(N__45654));
    LocalMux I__10628 (
            .O(N__45660),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    Odrv4 I__10627 (
            .O(N__45657),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    LocalMux I__10626 (
            .O(N__45654),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    InMux I__10625 (
            .O(N__45647),
            .I(N__45644));
    LocalMux I__10624 (
            .O(N__45644),
            .I(N__45641));
    Odrv12 I__10623 (
            .O(N__45641),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ));
    InMux I__10622 (
            .O(N__45638),
            .I(N__45632));
    InMux I__10621 (
            .O(N__45637),
            .I(N__45632));
    LocalMux I__10620 (
            .O(N__45632),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ));
    InMux I__10619 (
            .O(N__45629),
            .I(N__45623));
    InMux I__10618 (
            .O(N__45628),
            .I(N__45623));
    LocalMux I__10617 (
            .O(N__45623),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ));
    CascadeMux I__10616 (
            .O(N__45620),
            .I(N__45616));
    InMux I__10615 (
            .O(N__45619),
            .I(N__45610));
    InMux I__10614 (
            .O(N__45616),
            .I(N__45610));
    InMux I__10613 (
            .O(N__45615),
            .I(N__45607));
    LocalMux I__10612 (
            .O(N__45610),
            .I(N__45604));
    LocalMux I__10611 (
            .O(N__45607),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__10610 (
            .O(N__45604),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    CascadeMux I__10609 (
            .O(N__45599),
            .I(N__45595));
    InMux I__10608 (
            .O(N__45598),
            .I(N__45589));
    InMux I__10607 (
            .O(N__45595),
            .I(N__45589));
    InMux I__10606 (
            .O(N__45594),
            .I(N__45586));
    LocalMux I__10605 (
            .O(N__45589),
            .I(N__45583));
    LocalMux I__10604 (
            .O(N__45586),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__10603 (
            .O(N__45583),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    CascadeMux I__10602 (
            .O(N__45578),
            .I(N__45575));
    InMux I__10601 (
            .O(N__45575),
            .I(N__45572));
    LocalMux I__10600 (
            .O(N__45572),
            .I(N__45569));
    Odrv12 I__10599 (
            .O(N__45569),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt28 ));
    InMux I__10598 (
            .O(N__45566),
            .I(N__45563));
    LocalMux I__10597 (
            .O(N__45563),
            .I(N__45560));
    Odrv12 I__10596 (
            .O(N__45560),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt26 ));
    InMux I__10595 (
            .O(N__45557),
            .I(N__45552));
    InMux I__10594 (
            .O(N__45556),
            .I(N__45549));
    InMux I__10593 (
            .O(N__45555),
            .I(N__45546));
    LocalMux I__10592 (
            .O(N__45552),
            .I(N__45543));
    LocalMux I__10591 (
            .O(N__45549),
            .I(N__45540));
    LocalMux I__10590 (
            .O(N__45546),
            .I(N__45536));
    Span4Mux_h I__10589 (
            .O(N__45543),
            .I(N__45531));
    Span4Mux_v I__10588 (
            .O(N__45540),
            .I(N__45531));
    CascadeMux I__10587 (
            .O(N__45539),
            .I(N__45528));
    Sp12to4 I__10586 (
            .O(N__45536),
            .I(N__45525));
    Span4Mux_v I__10585 (
            .O(N__45531),
            .I(N__45522));
    InMux I__10584 (
            .O(N__45528),
            .I(N__45519));
    Span12Mux_v I__10583 (
            .O(N__45525),
            .I(N__45516));
    Span4Mux_h I__10582 (
            .O(N__45522),
            .I(N__45513));
    LocalMux I__10581 (
            .O(N__45519),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv12 I__10580 (
            .O(N__45516),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__10579 (
            .O(N__45513),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__10578 (
            .O(N__45506),
            .I(N__45503));
    InMux I__10577 (
            .O(N__45503),
            .I(N__45500));
    LocalMux I__10576 (
            .O(N__45500),
            .I(N__45494));
    InMux I__10575 (
            .O(N__45499),
            .I(N__45489));
    InMux I__10574 (
            .O(N__45498),
            .I(N__45489));
    InMux I__10573 (
            .O(N__45497),
            .I(N__45485));
    Span4Mux_h I__10572 (
            .O(N__45494),
            .I(N__45482));
    LocalMux I__10571 (
            .O(N__45489),
            .I(N__45479));
    InMux I__10570 (
            .O(N__45488),
            .I(N__45476));
    LocalMux I__10569 (
            .O(N__45485),
            .I(N__45473));
    Span4Mux_h I__10568 (
            .O(N__45482),
            .I(N__45470));
    Span4Mux_h I__10567 (
            .O(N__45479),
            .I(N__45467));
    LocalMux I__10566 (
            .O(N__45476),
            .I(N__45462));
    Span4Mux_h I__10565 (
            .O(N__45473),
            .I(N__45462));
    Span4Mux_v I__10564 (
            .O(N__45470),
            .I(N__45457));
    Span4Mux_v I__10563 (
            .O(N__45467),
            .I(N__45457));
    Span4Mux_v I__10562 (
            .O(N__45462),
            .I(N__45454));
    Odrv4 I__10561 (
            .O(N__45457),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__10560 (
            .O(N__45454),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    CascadeMux I__10559 (
            .O(N__45449),
            .I(N__45445));
    InMux I__10558 (
            .O(N__45448),
            .I(N__45440));
    InMux I__10557 (
            .O(N__45445),
            .I(N__45440));
    LocalMux I__10556 (
            .O(N__45440),
            .I(N__45437));
    Span4Mux_h I__10555 (
            .O(N__45437),
            .I(N__45433));
    InMux I__10554 (
            .O(N__45436),
            .I(N__45430));
    Span4Mux_h I__10553 (
            .O(N__45433),
            .I(N__45427));
    LocalMux I__10552 (
            .O(N__45430),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__10551 (
            .O(N__45427),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    CascadeMux I__10550 (
            .O(N__45422),
            .I(N__45419));
    InMux I__10549 (
            .O(N__45419),
            .I(N__45415));
    InMux I__10548 (
            .O(N__45418),
            .I(N__45412));
    LocalMux I__10547 (
            .O(N__45415),
            .I(N__45407));
    LocalMux I__10546 (
            .O(N__45412),
            .I(N__45407));
    Span4Mux_h I__10545 (
            .O(N__45407),
            .I(N__45403));
    InMux I__10544 (
            .O(N__45406),
            .I(N__45400));
    Span4Mux_h I__10543 (
            .O(N__45403),
            .I(N__45397));
    LocalMux I__10542 (
            .O(N__45400),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__10541 (
            .O(N__45397),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__10540 (
            .O(N__45392),
            .I(N__45389));
    LocalMux I__10539 (
            .O(N__45389),
            .I(N__45386));
    Span4Mux_h I__10538 (
            .O(N__45386),
            .I(N__45383));
    Odrv4 I__10537 (
            .O(N__45383),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ));
    InMux I__10536 (
            .O(N__45380),
            .I(N__45377));
    LocalMux I__10535 (
            .O(N__45377),
            .I(N__45374));
    Odrv12 I__10534 (
            .O(N__45374),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ));
    InMux I__10533 (
            .O(N__45371),
            .I(N__45365));
    InMux I__10532 (
            .O(N__45370),
            .I(N__45365));
    LocalMux I__10531 (
            .O(N__45365),
            .I(N__45362));
    Span4Mux_h I__10530 (
            .O(N__45362),
            .I(N__45358));
    InMux I__10529 (
            .O(N__45361),
            .I(N__45355));
    Span4Mux_h I__10528 (
            .O(N__45358),
            .I(N__45352));
    LocalMux I__10527 (
            .O(N__45355),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv4 I__10526 (
            .O(N__45352),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    CascadeMux I__10525 (
            .O(N__45347),
            .I(N__45343));
    InMux I__10524 (
            .O(N__45346),
            .I(N__45338));
    InMux I__10523 (
            .O(N__45343),
            .I(N__45338));
    LocalMux I__10522 (
            .O(N__45338),
            .I(N__45334));
    InMux I__10521 (
            .O(N__45337),
            .I(N__45331));
    Span12Mux_s10_v I__10520 (
            .O(N__45334),
            .I(N__45328));
    LocalMux I__10519 (
            .O(N__45331),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv12 I__10518 (
            .O(N__45328),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    CascadeMux I__10517 (
            .O(N__45323),
            .I(N__45320));
    InMux I__10516 (
            .O(N__45320),
            .I(N__45317));
    LocalMux I__10515 (
            .O(N__45317),
            .I(N__45314));
    Odrv12 I__10514 (
            .O(N__45314),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt26 ));
    InMux I__10513 (
            .O(N__45311),
            .I(N__45305));
    InMux I__10512 (
            .O(N__45310),
            .I(N__45305));
    LocalMux I__10511 (
            .O(N__45305),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ));
    InMux I__10510 (
            .O(N__45302),
            .I(N__45299));
    LocalMux I__10509 (
            .O(N__45299),
            .I(N__45296));
    Span4Mux_h I__10508 (
            .O(N__45296),
            .I(N__45293));
    Span4Mux_h I__10507 (
            .O(N__45293),
            .I(N__45290));
    Odrv4 I__10506 (
            .O(N__45290),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt28 ));
    InMux I__10505 (
            .O(N__45287),
            .I(N__45281));
    InMux I__10504 (
            .O(N__45286),
            .I(N__45281));
    LocalMux I__10503 (
            .O(N__45281),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    InMux I__10502 (
            .O(N__45278),
            .I(N__45273));
    InMux I__10501 (
            .O(N__45277),
            .I(N__45270));
    InMux I__10500 (
            .O(N__45276),
            .I(N__45267));
    LocalMux I__10499 (
            .O(N__45273),
            .I(N__45262));
    LocalMux I__10498 (
            .O(N__45270),
            .I(N__45262));
    LocalMux I__10497 (
            .O(N__45267),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv12 I__10496 (
            .O(N__45262),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    CascadeMux I__10495 (
            .O(N__45257),
            .I(N__45253));
    CascadeMux I__10494 (
            .O(N__45256),
            .I(N__45250));
    InMux I__10493 (
            .O(N__45253),
            .I(N__45247));
    InMux I__10492 (
            .O(N__45250),
            .I(N__45244));
    LocalMux I__10491 (
            .O(N__45247),
            .I(N__45238));
    LocalMux I__10490 (
            .O(N__45244),
            .I(N__45238));
    InMux I__10489 (
            .O(N__45243),
            .I(N__45235));
    Span4Mux_h I__10488 (
            .O(N__45238),
            .I(N__45232));
    LocalMux I__10487 (
            .O(N__45235),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__10486 (
            .O(N__45232),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__10485 (
            .O(N__45227),
            .I(N__45221));
    InMux I__10484 (
            .O(N__45226),
            .I(N__45221));
    LocalMux I__10483 (
            .O(N__45221),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    InMux I__10482 (
            .O(N__45218),
            .I(N__45212));
    InMux I__10481 (
            .O(N__45217),
            .I(N__45212));
    LocalMux I__10480 (
            .O(N__45212),
            .I(N__45208));
    InMux I__10479 (
            .O(N__45211),
            .I(N__45205));
    Span4Mux_v I__10478 (
            .O(N__45208),
            .I(N__45202));
    LocalMux I__10477 (
            .O(N__45205),
            .I(N__45199));
    Odrv4 I__10476 (
            .O(N__45202),
            .I(\current_shift_inst.un4_control_input1_2 ));
    Odrv12 I__10475 (
            .O(N__45199),
            .I(\current_shift_inst.un4_control_input1_2 ));
    InMux I__10474 (
            .O(N__45194),
            .I(N__45191));
    LocalMux I__10473 (
            .O(N__45191),
            .I(N__45187));
    CascadeMux I__10472 (
            .O(N__45190),
            .I(N__45183));
    Span4Mux_h I__10471 (
            .O(N__45187),
            .I(N__45179));
    InMux I__10470 (
            .O(N__45186),
            .I(N__45172));
    InMux I__10469 (
            .O(N__45183),
            .I(N__45172));
    InMux I__10468 (
            .O(N__45182),
            .I(N__45172));
    Odrv4 I__10467 (
            .O(N__45179),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__10466 (
            .O(N__45172),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__10465 (
            .O(N__45167),
            .I(N__45163));
    InMux I__10464 (
            .O(N__45166),
            .I(N__45158));
    InMux I__10463 (
            .O(N__45163),
            .I(N__45158));
    LocalMux I__10462 (
            .O(N__45158),
            .I(N__45154));
    InMux I__10461 (
            .O(N__45157),
            .I(N__45151));
    Span4Mux_v I__10460 (
            .O(N__45154),
            .I(N__45147));
    LocalMux I__10459 (
            .O(N__45151),
            .I(N__45144));
    InMux I__10458 (
            .O(N__45150),
            .I(N__45141));
    Span4Mux_h I__10457 (
            .O(N__45147),
            .I(N__45136));
    Span4Mux_h I__10456 (
            .O(N__45144),
            .I(N__45136));
    LocalMux I__10455 (
            .O(N__45141),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__10454 (
            .O(N__45136),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__10453 (
            .O(N__45131),
            .I(N__45128));
    InMux I__10452 (
            .O(N__45128),
            .I(N__45125));
    LocalMux I__10451 (
            .O(N__45125),
            .I(N__45122));
    Span4Mux_h I__10450 (
            .O(N__45122),
            .I(N__45119));
    Span4Mux_h I__10449 (
            .O(N__45119),
            .I(N__45116));
    Odrv4 I__10448 (
            .O(N__45116),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    CascadeMux I__10447 (
            .O(N__45113),
            .I(N__45110));
    InMux I__10446 (
            .O(N__45110),
            .I(N__45107));
    LocalMux I__10445 (
            .O(N__45107),
            .I(N__45104));
    Odrv12 I__10444 (
            .O(N__45104),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    InMux I__10443 (
            .O(N__45101),
            .I(N__45095));
    InMux I__10442 (
            .O(N__45100),
            .I(N__45095));
    LocalMux I__10441 (
            .O(N__45095),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    CascadeMux I__10440 (
            .O(N__45092),
            .I(N__45089));
    InMux I__10439 (
            .O(N__45089),
            .I(N__45083));
    InMux I__10438 (
            .O(N__45088),
            .I(N__45083));
    LocalMux I__10437 (
            .O(N__45083),
            .I(N__45080));
    Span4Mux_v I__10436 (
            .O(N__45080),
            .I(N__45076));
    InMux I__10435 (
            .O(N__45079),
            .I(N__45073));
    Sp12to4 I__10434 (
            .O(N__45076),
            .I(N__45066));
    LocalMux I__10433 (
            .O(N__45073),
            .I(N__45066));
    InMux I__10432 (
            .O(N__45072),
            .I(N__45061));
    InMux I__10431 (
            .O(N__45071),
            .I(N__45061));
    Odrv12 I__10430 (
            .O(N__45066),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__10429 (
            .O(N__45061),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__10428 (
            .O(N__45056),
            .I(N__45047));
    CascadeMux I__10427 (
            .O(N__45055),
            .I(N__45040));
    CascadeMux I__10426 (
            .O(N__45054),
            .I(N__45024));
    CascadeMux I__10425 (
            .O(N__45053),
            .I(N__45020));
    CascadeMux I__10424 (
            .O(N__45052),
            .I(N__45016));
    CascadeMux I__10423 (
            .O(N__45051),
            .I(N__45000));
    InMux I__10422 (
            .O(N__45050),
            .I(N__44989));
    InMux I__10421 (
            .O(N__45047),
            .I(N__44989));
    CascadeMux I__10420 (
            .O(N__45046),
            .I(N__44986));
    CascadeMux I__10419 (
            .O(N__45045),
            .I(N__44983));
    CascadeMux I__10418 (
            .O(N__45044),
            .I(N__44980));
    CascadeMux I__10417 (
            .O(N__45043),
            .I(N__44976));
    InMux I__10416 (
            .O(N__45040),
            .I(N__44966));
    CascadeMux I__10415 (
            .O(N__45039),
            .I(N__44962));
    CascadeMux I__10414 (
            .O(N__45038),
            .I(N__44958));
    CascadeMux I__10413 (
            .O(N__45037),
            .I(N__44955));
    InMux I__10412 (
            .O(N__45036),
            .I(N__44949));
    InMux I__10411 (
            .O(N__45035),
            .I(N__44949));
    InMux I__10410 (
            .O(N__45034),
            .I(N__44939));
    InMux I__10409 (
            .O(N__45033),
            .I(N__44939));
    InMux I__10408 (
            .O(N__45032),
            .I(N__44939));
    InMux I__10407 (
            .O(N__45031),
            .I(N__44939));
    CascadeMux I__10406 (
            .O(N__45030),
            .I(N__44928));
    CascadeMux I__10405 (
            .O(N__45029),
            .I(N__44920));
    InMux I__10404 (
            .O(N__45028),
            .I(N__44902));
    InMux I__10403 (
            .O(N__45027),
            .I(N__44902));
    InMux I__10402 (
            .O(N__45024),
            .I(N__44902));
    InMux I__10401 (
            .O(N__45023),
            .I(N__44902));
    InMux I__10400 (
            .O(N__45020),
            .I(N__44902));
    InMux I__10399 (
            .O(N__45019),
            .I(N__44902));
    InMux I__10398 (
            .O(N__45016),
            .I(N__44902));
    InMux I__10397 (
            .O(N__45015),
            .I(N__44902));
    CascadeMux I__10396 (
            .O(N__45014),
            .I(N__44899));
    CascadeMux I__10395 (
            .O(N__45013),
            .I(N__44895));
    CascadeMux I__10394 (
            .O(N__45012),
            .I(N__44891));
    CascadeMux I__10393 (
            .O(N__45011),
            .I(N__44887));
    CascadeMux I__10392 (
            .O(N__45010),
            .I(N__44883));
    CascadeMux I__10391 (
            .O(N__45009),
            .I(N__44879));
    CascadeMux I__10390 (
            .O(N__45008),
            .I(N__44875));
    CascadeMux I__10389 (
            .O(N__45007),
            .I(N__44871));
    CascadeMux I__10388 (
            .O(N__45006),
            .I(N__44867));
    CascadeMux I__10387 (
            .O(N__45005),
            .I(N__44863));
    CascadeMux I__10386 (
            .O(N__45004),
            .I(N__44859));
    InMux I__10385 (
            .O(N__45003),
            .I(N__44853));
    InMux I__10384 (
            .O(N__45000),
            .I(N__44853));
    CascadeMux I__10383 (
            .O(N__44999),
            .I(N__44847));
    CascadeMux I__10382 (
            .O(N__44998),
            .I(N__44844));
    CascadeMux I__10381 (
            .O(N__44997),
            .I(N__44841));
    CascadeMux I__10380 (
            .O(N__44996),
            .I(N__44838));
    CascadeMux I__10379 (
            .O(N__44995),
            .I(N__44835));
    CascadeMux I__10378 (
            .O(N__44994),
            .I(N__44830));
    LocalMux I__10377 (
            .O(N__44989),
            .I(N__44824));
    InMux I__10376 (
            .O(N__44986),
            .I(N__44821));
    InMux I__10375 (
            .O(N__44983),
            .I(N__44818));
    InMux I__10374 (
            .O(N__44980),
            .I(N__44811));
    InMux I__10373 (
            .O(N__44979),
            .I(N__44811));
    InMux I__10372 (
            .O(N__44976),
            .I(N__44811));
    CascadeMux I__10371 (
            .O(N__44975),
            .I(N__44807));
    CascadeMux I__10370 (
            .O(N__44974),
            .I(N__44803));
    CascadeMux I__10369 (
            .O(N__44973),
            .I(N__44799));
    CascadeMux I__10368 (
            .O(N__44972),
            .I(N__44795));
    CascadeMux I__10367 (
            .O(N__44971),
            .I(N__44791));
    CascadeMux I__10366 (
            .O(N__44970),
            .I(N__44787));
    CascadeMux I__10365 (
            .O(N__44969),
            .I(N__44783));
    LocalMux I__10364 (
            .O(N__44966),
            .I(N__44772));
    InMux I__10363 (
            .O(N__44965),
            .I(N__44769));
    InMux I__10362 (
            .O(N__44962),
            .I(N__44764));
    InMux I__10361 (
            .O(N__44961),
            .I(N__44764));
    InMux I__10360 (
            .O(N__44958),
            .I(N__44761));
    InMux I__10359 (
            .O(N__44955),
            .I(N__44756));
    InMux I__10358 (
            .O(N__44954),
            .I(N__44756));
    LocalMux I__10357 (
            .O(N__44949),
            .I(N__44753));
    InMux I__10356 (
            .O(N__44948),
            .I(N__44750));
    LocalMux I__10355 (
            .O(N__44939),
            .I(N__44747));
    InMux I__10354 (
            .O(N__44938),
            .I(N__44732));
    InMux I__10353 (
            .O(N__44937),
            .I(N__44732));
    InMux I__10352 (
            .O(N__44936),
            .I(N__44732));
    InMux I__10351 (
            .O(N__44935),
            .I(N__44732));
    InMux I__10350 (
            .O(N__44934),
            .I(N__44732));
    InMux I__10349 (
            .O(N__44933),
            .I(N__44732));
    InMux I__10348 (
            .O(N__44932),
            .I(N__44732));
    InMux I__10347 (
            .O(N__44931),
            .I(N__44717));
    InMux I__10346 (
            .O(N__44928),
            .I(N__44717));
    InMux I__10345 (
            .O(N__44927),
            .I(N__44717));
    InMux I__10344 (
            .O(N__44926),
            .I(N__44717));
    InMux I__10343 (
            .O(N__44925),
            .I(N__44717));
    InMux I__10342 (
            .O(N__44924),
            .I(N__44717));
    InMux I__10341 (
            .O(N__44923),
            .I(N__44717));
    InMux I__10340 (
            .O(N__44920),
            .I(N__44712));
    InMux I__10339 (
            .O(N__44919),
            .I(N__44712));
    LocalMux I__10338 (
            .O(N__44902),
            .I(N__44709));
    InMux I__10337 (
            .O(N__44899),
            .I(N__44692));
    InMux I__10336 (
            .O(N__44898),
            .I(N__44692));
    InMux I__10335 (
            .O(N__44895),
            .I(N__44692));
    InMux I__10334 (
            .O(N__44894),
            .I(N__44692));
    InMux I__10333 (
            .O(N__44891),
            .I(N__44692));
    InMux I__10332 (
            .O(N__44890),
            .I(N__44692));
    InMux I__10331 (
            .O(N__44887),
            .I(N__44692));
    InMux I__10330 (
            .O(N__44886),
            .I(N__44692));
    InMux I__10329 (
            .O(N__44883),
            .I(N__44675));
    InMux I__10328 (
            .O(N__44882),
            .I(N__44675));
    InMux I__10327 (
            .O(N__44879),
            .I(N__44675));
    InMux I__10326 (
            .O(N__44878),
            .I(N__44675));
    InMux I__10325 (
            .O(N__44875),
            .I(N__44675));
    InMux I__10324 (
            .O(N__44874),
            .I(N__44675));
    InMux I__10323 (
            .O(N__44871),
            .I(N__44675));
    InMux I__10322 (
            .O(N__44870),
            .I(N__44675));
    InMux I__10321 (
            .O(N__44867),
            .I(N__44662));
    InMux I__10320 (
            .O(N__44866),
            .I(N__44662));
    InMux I__10319 (
            .O(N__44863),
            .I(N__44662));
    InMux I__10318 (
            .O(N__44862),
            .I(N__44662));
    InMux I__10317 (
            .O(N__44859),
            .I(N__44662));
    InMux I__10316 (
            .O(N__44858),
            .I(N__44662));
    LocalMux I__10315 (
            .O(N__44853),
            .I(N__44659));
    InMux I__10314 (
            .O(N__44852),
            .I(N__44652));
    InMux I__10313 (
            .O(N__44851),
            .I(N__44652));
    InMux I__10312 (
            .O(N__44850),
            .I(N__44652));
    InMux I__10311 (
            .O(N__44847),
            .I(N__44645));
    InMux I__10310 (
            .O(N__44844),
            .I(N__44645));
    InMux I__10309 (
            .O(N__44841),
            .I(N__44645));
    InMux I__10308 (
            .O(N__44838),
            .I(N__44628));
    InMux I__10307 (
            .O(N__44835),
            .I(N__44628));
    InMux I__10306 (
            .O(N__44834),
            .I(N__44628));
    InMux I__10305 (
            .O(N__44833),
            .I(N__44628));
    InMux I__10304 (
            .O(N__44830),
            .I(N__44628));
    InMux I__10303 (
            .O(N__44829),
            .I(N__44628));
    InMux I__10302 (
            .O(N__44828),
            .I(N__44628));
    InMux I__10301 (
            .O(N__44827),
            .I(N__44628));
    Span4Mux_v I__10300 (
            .O(N__44824),
            .I(N__44619));
    LocalMux I__10299 (
            .O(N__44821),
            .I(N__44612));
    LocalMux I__10298 (
            .O(N__44818),
            .I(N__44612));
    LocalMux I__10297 (
            .O(N__44811),
            .I(N__44612));
    InMux I__10296 (
            .O(N__44810),
            .I(N__44597));
    InMux I__10295 (
            .O(N__44807),
            .I(N__44597));
    InMux I__10294 (
            .O(N__44806),
            .I(N__44597));
    InMux I__10293 (
            .O(N__44803),
            .I(N__44597));
    InMux I__10292 (
            .O(N__44802),
            .I(N__44597));
    InMux I__10291 (
            .O(N__44799),
            .I(N__44597));
    InMux I__10290 (
            .O(N__44798),
            .I(N__44597));
    InMux I__10289 (
            .O(N__44795),
            .I(N__44580));
    InMux I__10288 (
            .O(N__44794),
            .I(N__44580));
    InMux I__10287 (
            .O(N__44791),
            .I(N__44580));
    InMux I__10286 (
            .O(N__44790),
            .I(N__44580));
    InMux I__10285 (
            .O(N__44787),
            .I(N__44580));
    InMux I__10284 (
            .O(N__44786),
            .I(N__44580));
    InMux I__10283 (
            .O(N__44783),
            .I(N__44580));
    InMux I__10282 (
            .O(N__44782),
            .I(N__44580));
    CascadeMux I__10281 (
            .O(N__44781),
            .I(N__44577));
    CascadeMux I__10280 (
            .O(N__44780),
            .I(N__44573));
    CascadeMux I__10279 (
            .O(N__44779),
            .I(N__44569));
    CascadeMux I__10278 (
            .O(N__44778),
            .I(N__44565));
    CascadeMux I__10277 (
            .O(N__44777),
            .I(N__44561));
    CascadeMux I__10276 (
            .O(N__44776),
            .I(N__44557));
    CascadeMux I__10275 (
            .O(N__44775),
            .I(N__44553));
    Span4Mux_h I__10274 (
            .O(N__44772),
            .I(N__44545));
    LocalMux I__10273 (
            .O(N__44769),
            .I(N__44545));
    LocalMux I__10272 (
            .O(N__44764),
            .I(N__44545));
    LocalMux I__10271 (
            .O(N__44761),
            .I(N__44542));
    LocalMux I__10270 (
            .O(N__44756),
            .I(N__44539));
    Span4Mux_h I__10269 (
            .O(N__44753),
            .I(N__44518));
    LocalMux I__10268 (
            .O(N__44750),
            .I(N__44518));
    Span4Mux_h I__10267 (
            .O(N__44747),
            .I(N__44518));
    LocalMux I__10266 (
            .O(N__44732),
            .I(N__44518));
    LocalMux I__10265 (
            .O(N__44717),
            .I(N__44518));
    LocalMux I__10264 (
            .O(N__44712),
            .I(N__44518));
    Span4Mux_v I__10263 (
            .O(N__44709),
            .I(N__44518));
    LocalMux I__10262 (
            .O(N__44692),
            .I(N__44518));
    LocalMux I__10261 (
            .O(N__44675),
            .I(N__44518));
    LocalMux I__10260 (
            .O(N__44662),
            .I(N__44518));
    Span4Mux_h I__10259 (
            .O(N__44659),
            .I(N__44515));
    LocalMux I__10258 (
            .O(N__44652),
            .I(N__44508));
    LocalMux I__10257 (
            .O(N__44645),
            .I(N__44508));
    LocalMux I__10256 (
            .O(N__44628),
            .I(N__44508));
    InMux I__10255 (
            .O(N__44627),
            .I(N__44505));
    InMux I__10254 (
            .O(N__44626),
            .I(N__44494));
    InMux I__10253 (
            .O(N__44625),
            .I(N__44494));
    InMux I__10252 (
            .O(N__44624),
            .I(N__44494));
    InMux I__10251 (
            .O(N__44623),
            .I(N__44494));
    InMux I__10250 (
            .O(N__44622),
            .I(N__44494));
    Span4Mux_h I__10249 (
            .O(N__44619),
            .I(N__44485));
    Span4Mux_v I__10248 (
            .O(N__44612),
            .I(N__44485));
    LocalMux I__10247 (
            .O(N__44597),
            .I(N__44485));
    LocalMux I__10246 (
            .O(N__44580),
            .I(N__44485));
    InMux I__10245 (
            .O(N__44577),
            .I(N__44468));
    InMux I__10244 (
            .O(N__44576),
            .I(N__44468));
    InMux I__10243 (
            .O(N__44573),
            .I(N__44468));
    InMux I__10242 (
            .O(N__44572),
            .I(N__44468));
    InMux I__10241 (
            .O(N__44569),
            .I(N__44468));
    InMux I__10240 (
            .O(N__44568),
            .I(N__44468));
    InMux I__10239 (
            .O(N__44565),
            .I(N__44468));
    InMux I__10238 (
            .O(N__44564),
            .I(N__44468));
    InMux I__10237 (
            .O(N__44561),
            .I(N__44455));
    InMux I__10236 (
            .O(N__44560),
            .I(N__44455));
    InMux I__10235 (
            .O(N__44557),
            .I(N__44455));
    InMux I__10234 (
            .O(N__44556),
            .I(N__44455));
    InMux I__10233 (
            .O(N__44553),
            .I(N__44455));
    InMux I__10232 (
            .O(N__44552),
            .I(N__44455));
    Span4Mux_v I__10231 (
            .O(N__44545),
            .I(N__44446));
    Span4Mux_v I__10230 (
            .O(N__44542),
            .I(N__44446));
    Span4Mux_h I__10229 (
            .O(N__44539),
            .I(N__44446));
    Span4Mux_v I__10228 (
            .O(N__44518),
            .I(N__44446));
    Odrv4 I__10227 (
            .O(N__44515),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10226 (
            .O(N__44508),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10225 (
            .O(N__44505),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10224 (
            .O(N__44494),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10223 (
            .O(N__44485),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10222 (
            .O(N__44468),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__10221 (
            .O(N__44455),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__10220 (
            .O(N__44446),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__10219 (
            .O(N__44429),
            .I(N__44411));
    CascadeMux I__10218 (
            .O(N__44428),
            .I(N__44408));
    InMux I__10217 (
            .O(N__44427),
            .I(N__44385));
    InMux I__10216 (
            .O(N__44426),
            .I(N__44382));
    InMux I__10215 (
            .O(N__44425),
            .I(N__44369));
    InMux I__10214 (
            .O(N__44424),
            .I(N__44369));
    InMux I__10213 (
            .O(N__44423),
            .I(N__44369));
    InMux I__10212 (
            .O(N__44422),
            .I(N__44369));
    InMux I__10211 (
            .O(N__44421),
            .I(N__44369));
    InMux I__10210 (
            .O(N__44420),
            .I(N__44369));
    CascadeMux I__10209 (
            .O(N__44419),
            .I(N__44366));
    InMux I__10208 (
            .O(N__44418),
            .I(N__44356));
    InMux I__10207 (
            .O(N__44417),
            .I(N__44352));
    CascadeMux I__10206 (
            .O(N__44416),
            .I(N__44349));
    InMux I__10205 (
            .O(N__44415),
            .I(N__44344));
    InMux I__10204 (
            .O(N__44414),
            .I(N__44344));
    InMux I__10203 (
            .O(N__44411),
            .I(N__44339));
    InMux I__10202 (
            .O(N__44408),
            .I(N__44339));
    InMux I__10201 (
            .O(N__44407),
            .I(N__44336));
    InMux I__10200 (
            .O(N__44406),
            .I(N__44323));
    InMux I__10199 (
            .O(N__44405),
            .I(N__44323));
    InMux I__10198 (
            .O(N__44404),
            .I(N__44323));
    InMux I__10197 (
            .O(N__44403),
            .I(N__44323));
    InMux I__10196 (
            .O(N__44402),
            .I(N__44323));
    InMux I__10195 (
            .O(N__44401),
            .I(N__44323));
    InMux I__10194 (
            .O(N__44400),
            .I(N__44316));
    InMux I__10193 (
            .O(N__44399),
            .I(N__44316));
    InMux I__10192 (
            .O(N__44398),
            .I(N__44316));
    InMux I__10191 (
            .O(N__44397),
            .I(N__44311));
    InMux I__10190 (
            .O(N__44396),
            .I(N__44311));
    InMux I__10189 (
            .O(N__44395),
            .I(N__44302));
    InMux I__10188 (
            .O(N__44394),
            .I(N__44302));
    InMux I__10187 (
            .O(N__44393),
            .I(N__44302));
    InMux I__10186 (
            .O(N__44392),
            .I(N__44302));
    InMux I__10185 (
            .O(N__44391),
            .I(N__44299));
    InMux I__10184 (
            .O(N__44390),
            .I(N__44288));
    InMux I__10183 (
            .O(N__44389),
            .I(N__44283));
    InMux I__10182 (
            .O(N__44388),
            .I(N__44283));
    LocalMux I__10181 (
            .O(N__44385),
            .I(N__44272));
    LocalMux I__10180 (
            .O(N__44382),
            .I(N__44272));
    LocalMux I__10179 (
            .O(N__44369),
            .I(N__44269));
    InMux I__10178 (
            .O(N__44366),
            .I(N__44252));
    InMux I__10177 (
            .O(N__44365),
            .I(N__44252));
    InMux I__10176 (
            .O(N__44364),
            .I(N__44252));
    InMux I__10175 (
            .O(N__44363),
            .I(N__44252));
    InMux I__10174 (
            .O(N__44362),
            .I(N__44252));
    InMux I__10173 (
            .O(N__44361),
            .I(N__44252));
    InMux I__10172 (
            .O(N__44360),
            .I(N__44252));
    InMux I__10171 (
            .O(N__44359),
            .I(N__44252));
    LocalMux I__10170 (
            .O(N__44356),
            .I(N__44249));
    InMux I__10169 (
            .O(N__44355),
            .I(N__44246));
    LocalMux I__10168 (
            .O(N__44352),
            .I(N__44243));
    InMux I__10167 (
            .O(N__44349),
            .I(N__44240));
    LocalMux I__10166 (
            .O(N__44344),
            .I(N__44236));
    LocalMux I__10165 (
            .O(N__44339),
            .I(N__44227));
    LocalMux I__10164 (
            .O(N__44336),
            .I(N__44227));
    LocalMux I__10163 (
            .O(N__44323),
            .I(N__44227));
    LocalMux I__10162 (
            .O(N__44316),
            .I(N__44227));
    LocalMux I__10161 (
            .O(N__44311),
            .I(N__44222));
    LocalMux I__10160 (
            .O(N__44302),
            .I(N__44222));
    LocalMux I__10159 (
            .O(N__44299),
            .I(N__44219));
    InMux I__10158 (
            .O(N__44298),
            .I(N__44216));
    InMux I__10157 (
            .O(N__44297),
            .I(N__44201));
    InMux I__10156 (
            .O(N__44296),
            .I(N__44201));
    InMux I__10155 (
            .O(N__44295),
            .I(N__44201));
    InMux I__10154 (
            .O(N__44294),
            .I(N__44201));
    InMux I__10153 (
            .O(N__44293),
            .I(N__44201));
    InMux I__10152 (
            .O(N__44292),
            .I(N__44201));
    InMux I__10151 (
            .O(N__44291),
            .I(N__44201));
    LocalMux I__10150 (
            .O(N__44288),
            .I(N__44184));
    LocalMux I__10149 (
            .O(N__44283),
            .I(N__44184));
    InMux I__10148 (
            .O(N__44282),
            .I(N__44171));
    InMux I__10147 (
            .O(N__44281),
            .I(N__44171));
    InMux I__10146 (
            .O(N__44280),
            .I(N__44171));
    InMux I__10145 (
            .O(N__44279),
            .I(N__44171));
    InMux I__10144 (
            .O(N__44278),
            .I(N__44171));
    InMux I__10143 (
            .O(N__44277),
            .I(N__44171));
    Span4Mux_v I__10142 (
            .O(N__44272),
            .I(N__44162));
    Span4Mux_v I__10141 (
            .O(N__44269),
            .I(N__44162));
    LocalMux I__10140 (
            .O(N__44252),
            .I(N__44162));
    Span4Mux_h I__10139 (
            .O(N__44249),
            .I(N__44162));
    LocalMux I__10138 (
            .O(N__44246),
            .I(N__44155));
    Span4Mux_h I__10137 (
            .O(N__44243),
            .I(N__44155));
    LocalMux I__10136 (
            .O(N__44240),
            .I(N__44155));
    InMux I__10135 (
            .O(N__44239),
            .I(N__44152));
    Span4Mux_v I__10134 (
            .O(N__44236),
            .I(N__44145));
    Span4Mux_v I__10133 (
            .O(N__44227),
            .I(N__44145));
    Span4Mux_v I__10132 (
            .O(N__44222),
            .I(N__44145));
    Span4Mux_v I__10131 (
            .O(N__44219),
            .I(N__44138));
    LocalMux I__10130 (
            .O(N__44216),
            .I(N__44138));
    LocalMux I__10129 (
            .O(N__44201),
            .I(N__44138));
    InMux I__10128 (
            .O(N__44200),
            .I(N__44123));
    InMux I__10127 (
            .O(N__44199),
            .I(N__44123));
    InMux I__10126 (
            .O(N__44198),
            .I(N__44123));
    InMux I__10125 (
            .O(N__44197),
            .I(N__44123));
    InMux I__10124 (
            .O(N__44196),
            .I(N__44123));
    InMux I__10123 (
            .O(N__44195),
            .I(N__44123));
    InMux I__10122 (
            .O(N__44194),
            .I(N__44123));
    InMux I__10121 (
            .O(N__44193),
            .I(N__44118));
    InMux I__10120 (
            .O(N__44192),
            .I(N__44118));
    InMux I__10119 (
            .O(N__44191),
            .I(N__44115));
    InMux I__10118 (
            .O(N__44190),
            .I(N__44110));
    InMux I__10117 (
            .O(N__44189),
            .I(N__44110));
    Span4Mux_v I__10116 (
            .O(N__44184),
            .I(N__44105));
    LocalMux I__10115 (
            .O(N__44171),
            .I(N__44105));
    Span4Mux_h I__10114 (
            .O(N__44162),
            .I(N__44102));
    Span4Mux_v I__10113 (
            .O(N__44155),
            .I(N__44095));
    LocalMux I__10112 (
            .O(N__44152),
            .I(N__44095));
    Span4Mux_h I__10111 (
            .O(N__44145),
            .I(N__44095));
    Odrv4 I__10110 (
            .O(N__44138),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10109 (
            .O(N__44123),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10108 (
            .O(N__44118),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10107 (
            .O(N__44115),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10106 (
            .O(N__44110),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10105 (
            .O(N__44105),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10104 (
            .O(N__44102),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10103 (
            .O(N__44095),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__10102 (
            .O(N__44078),
            .I(N__44075));
    InMux I__10101 (
            .O(N__44075),
            .I(N__44072));
    LocalMux I__10100 (
            .O(N__44072),
            .I(N__44069));
    Span4Mux_h I__10099 (
            .O(N__44069),
            .I(N__44066));
    Odrv4 I__10098 (
            .O(N__44066),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__10097 (
            .O(N__44063),
            .I(N__44058));
    InMux I__10096 (
            .O(N__44062),
            .I(N__44055));
    InMux I__10095 (
            .O(N__44061),
            .I(N__44052));
    LocalMux I__10094 (
            .O(N__44058),
            .I(N__44047));
    LocalMux I__10093 (
            .O(N__44055),
            .I(N__44047));
    LocalMux I__10092 (
            .O(N__44052),
            .I(N__44043));
    Span4Mux_h I__10091 (
            .O(N__44047),
            .I(N__44040));
    InMux I__10090 (
            .O(N__44046),
            .I(N__44037));
    Span4Mux_v I__10089 (
            .O(N__44043),
            .I(N__44034));
    Span4Mux_v I__10088 (
            .O(N__44040),
            .I(N__44029));
    LocalMux I__10087 (
            .O(N__44037),
            .I(N__44029));
    Odrv4 I__10086 (
            .O(N__44034),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    Odrv4 I__10085 (
            .O(N__44029),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__10084 (
            .O(N__44024),
            .I(N__44021));
    LocalMux I__10083 (
            .O(N__44021),
            .I(N__44018));
    Span4Mux_h I__10082 (
            .O(N__44018),
            .I(N__44015));
    Odrv4 I__10081 (
            .O(N__44015),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__10080 (
            .O(N__44012),
            .I(N__44009));
    LocalMux I__10079 (
            .O(N__44009),
            .I(N__44004));
    InMux I__10078 (
            .O(N__44008),
            .I(N__44001));
    InMux I__10077 (
            .O(N__44007),
            .I(N__43998));
    Span4Mux_h I__10076 (
            .O(N__44004),
            .I(N__43990));
    LocalMux I__10075 (
            .O(N__44001),
            .I(N__43990));
    LocalMux I__10074 (
            .O(N__43998),
            .I(N__43990));
    InMux I__10073 (
            .O(N__43997),
            .I(N__43987));
    Span4Mux_h I__10072 (
            .O(N__43990),
            .I(N__43982));
    LocalMux I__10071 (
            .O(N__43987),
            .I(N__43982));
    Span4Mux_v I__10070 (
            .O(N__43982),
            .I(N__43979));
    Odrv4 I__10069 (
            .O(N__43979),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__10068 (
            .O(N__43976),
            .I(N__43973));
    LocalMux I__10067 (
            .O(N__43973),
            .I(N__43970));
    Odrv4 I__10066 (
            .O(N__43970),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    CascadeMux I__10065 (
            .O(N__43967),
            .I(N__43963));
    CascadeMux I__10064 (
            .O(N__43966),
            .I(N__43960));
    InMux I__10063 (
            .O(N__43963),
            .I(N__43956));
    InMux I__10062 (
            .O(N__43960),
            .I(N__43953));
    InMux I__10061 (
            .O(N__43959),
            .I(N__43950));
    LocalMux I__10060 (
            .O(N__43956),
            .I(N__43946));
    LocalMux I__10059 (
            .O(N__43953),
            .I(N__43943));
    LocalMux I__10058 (
            .O(N__43950),
            .I(N__43940));
    InMux I__10057 (
            .O(N__43949),
            .I(N__43937));
    Span4Mux_h I__10056 (
            .O(N__43946),
            .I(N__43934));
    Span4Mux_v I__10055 (
            .O(N__43943),
            .I(N__43931));
    Span4Mux_h I__10054 (
            .O(N__43940),
            .I(N__43928));
    LocalMux I__10053 (
            .O(N__43937),
            .I(N__43925));
    Odrv4 I__10052 (
            .O(N__43934),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__10051 (
            .O(N__43931),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__10050 (
            .O(N__43928),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv12 I__10049 (
            .O(N__43925),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__10048 (
            .O(N__43916),
            .I(N__43913));
    LocalMux I__10047 (
            .O(N__43913),
            .I(N__43910));
    Odrv12 I__10046 (
            .O(N__43910),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    CascadeMux I__10045 (
            .O(N__43907),
            .I(N__43904));
    InMux I__10044 (
            .O(N__43904),
            .I(N__43901));
    LocalMux I__10043 (
            .O(N__43901),
            .I(N__43896));
    InMux I__10042 (
            .O(N__43900),
            .I(N__43891));
    InMux I__10041 (
            .O(N__43899),
            .I(N__43891));
    Span4Mux_h I__10040 (
            .O(N__43896),
            .I(N__43885));
    LocalMux I__10039 (
            .O(N__43891),
            .I(N__43885));
    InMux I__10038 (
            .O(N__43890),
            .I(N__43882));
    Span4Mux_h I__10037 (
            .O(N__43885),
            .I(N__43879));
    LocalMux I__10036 (
            .O(N__43882),
            .I(N__43876));
    Odrv4 I__10035 (
            .O(N__43879),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__10034 (
            .O(N__43876),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__10033 (
            .O(N__43871),
            .I(N__43868));
    LocalMux I__10032 (
            .O(N__43868),
            .I(N__43865));
    Odrv12 I__10031 (
            .O(N__43865),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__10030 (
            .O(N__43862),
            .I(N__43859));
    LocalMux I__10029 (
            .O(N__43859),
            .I(N__43856));
    Span4Mux_v I__10028 (
            .O(N__43856),
            .I(N__43852));
    CascadeMux I__10027 (
            .O(N__43855),
            .I(N__43848));
    Span4Mux_h I__10026 (
            .O(N__43852),
            .I(N__43840));
    InMux I__10025 (
            .O(N__43851),
            .I(N__43837));
    InMux I__10024 (
            .O(N__43848),
            .I(N__43830));
    InMux I__10023 (
            .O(N__43847),
            .I(N__43830));
    InMux I__10022 (
            .O(N__43846),
            .I(N__43830));
    InMux I__10021 (
            .O(N__43845),
            .I(N__43827));
    InMux I__10020 (
            .O(N__43844),
            .I(N__43822));
    InMux I__10019 (
            .O(N__43843),
            .I(N__43822));
    Span4Mux_h I__10018 (
            .O(N__43840),
            .I(N__43818));
    LocalMux I__10017 (
            .O(N__43837),
            .I(N__43811));
    LocalMux I__10016 (
            .O(N__43830),
            .I(N__43811));
    LocalMux I__10015 (
            .O(N__43827),
            .I(N__43811));
    LocalMux I__10014 (
            .O(N__43822),
            .I(N__43808));
    InMux I__10013 (
            .O(N__43821),
            .I(N__43805));
    Span4Mux_h I__10012 (
            .O(N__43818),
            .I(N__43799));
    Span4Mux_v I__10011 (
            .O(N__43811),
            .I(N__43799));
    Span4Mux_h I__10010 (
            .O(N__43808),
            .I(N__43796));
    LocalMux I__10009 (
            .O(N__43805),
            .I(N__43793));
    InMux I__10008 (
            .O(N__43804),
            .I(N__43790));
    Odrv4 I__10007 (
            .O(N__43799),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__10006 (
            .O(N__43796),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__10005 (
            .O(N__43793),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    LocalMux I__10004 (
            .O(N__43790),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    CascadeMux I__10003 (
            .O(N__43781),
            .I(N__43778));
    InMux I__10002 (
            .O(N__43778),
            .I(N__43775));
    LocalMux I__10001 (
            .O(N__43775),
            .I(N__43772));
    Span4Mux_h I__10000 (
            .O(N__43772),
            .I(N__43769));
    Odrv4 I__9999 (
            .O(N__43769),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt24 ));
    InMux I__9998 (
            .O(N__43766),
            .I(N__43763));
    LocalMux I__9997 (
            .O(N__43763),
            .I(N__43760));
    Span12Mux_v I__9996 (
            .O(N__43760),
            .I(N__43757));
    Odrv12 I__9995 (
            .O(N__43757),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    CascadeMux I__9994 (
            .O(N__43754),
            .I(N__43751));
    InMux I__9993 (
            .O(N__43751),
            .I(N__43747));
    CascadeMux I__9992 (
            .O(N__43750),
            .I(N__43744));
    LocalMux I__9991 (
            .O(N__43747),
            .I(N__43740));
    InMux I__9990 (
            .O(N__43744),
            .I(N__43735));
    InMux I__9989 (
            .O(N__43743),
            .I(N__43735));
    Odrv4 I__9988 (
            .O(N__43740),
            .I(\current_shift_inst.un4_control_input1_29 ));
    LocalMux I__9987 (
            .O(N__43735),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__9986 (
            .O(N__43730),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    CascadeMux I__9985 (
            .O(N__43727),
            .I(N__43723));
    InMux I__9984 (
            .O(N__43726),
            .I(N__43720));
    InMux I__9983 (
            .O(N__43723),
            .I(N__43717));
    LocalMux I__9982 (
            .O(N__43720),
            .I(N__43711));
    LocalMux I__9981 (
            .O(N__43717),
            .I(N__43711));
    InMux I__9980 (
            .O(N__43716),
            .I(N__43708));
    Odrv12 I__9979 (
            .O(N__43711),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__9978 (
            .O(N__43708),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__9977 (
            .O(N__43703),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__9976 (
            .O(N__43700),
            .I(\current_shift_inst.un4_control_input1_31 ));
    CascadeMux I__9975 (
            .O(N__43697),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ));
    InMux I__9974 (
            .O(N__43694),
            .I(N__43691));
    LocalMux I__9973 (
            .O(N__43691),
            .I(N__43688));
    Odrv4 I__9972 (
            .O(N__43688),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__9971 (
            .O(N__43685),
            .I(N__43681));
    InMux I__9970 (
            .O(N__43684),
            .I(N__43676));
    LocalMux I__9969 (
            .O(N__43681),
            .I(N__43673));
    InMux I__9968 (
            .O(N__43680),
            .I(N__43668));
    InMux I__9967 (
            .O(N__43679),
            .I(N__43668));
    LocalMux I__9966 (
            .O(N__43676),
            .I(N__43665));
    Span4Mux_h I__9965 (
            .O(N__43673),
            .I(N__43660));
    LocalMux I__9964 (
            .O(N__43668),
            .I(N__43660));
    Span4Mux_h I__9963 (
            .O(N__43665),
            .I(N__43657));
    Span4Mux_v I__9962 (
            .O(N__43660),
            .I(N__43654));
    Odrv4 I__9961 (
            .O(N__43657),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__9960 (
            .O(N__43654),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__9959 (
            .O(N__43649),
            .I(N__43646));
    LocalMux I__9958 (
            .O(N__43646),
            .I(N__43641));
    InMux I__9957 (
            .O(N__43645),
            .I(N__43638));
    InMux I__9956 (
            .O(N__43644),
            .I(N__43635));
    Odrv4 I__9955 (
            .O(N__43641),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__9954 (
            .O(N__43638),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__9953 (
            .O(N__43635),
            .I(\current_shift_inst.un4_control_input1_7 ));
    CascadeMux I__9952 (
            .O(N__43628),
            .I(N__43625));
    InMux I__9951 (
            .O(N__43625),
            .I(N__43622));
    LocalMux I__9950 (
            .O(N__43622),
            .I(N__43619));
    Span4Mux_h I__9949 (
            .O(N__43619),
            .I(N__43616));
    Span4Mux_v I__9948 (
            .O(N__43616),
            .I(N__43613));
    Odrv4 I__9947 (
            .O(N__43613),
            .I(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ));
    CascadeMux I__9946 (
            .O(N__43610),
            .I(N__43607));
    InMux I__9945 (
            .O(N__43607),
            .I(N__43604));
    LocalMux I__9944 (
            .O(N__43604),
            .I(N__43601));
    Span12Mux_v I__9943 (
            .O(N__43601),
            .I(N__43598));
    Odrv12 I__9942 (
            .O(N__43598),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ));
    InMux I__9941 (
            .O(N__43595),
            .I(N__43590));
    InMux I__9940 (
            .O(N__43594),
            .I(N__43587));
    InMux I__9939 (
            .O(N__43593),
            .I(N__43584));
    LocalMux I__9938 (
            .O(N__43590),
            .I(N__43581));
    LocalMux I__9937 (
            .O(N__43587),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__9936 (
            .O(N__43584),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv4 I__9935 (
            .O(N__43581),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    CEMux I__9934 (
            .O(N__43574),
            .I(N__43550));
    CEMux I__9933 (
            .O(N__43573),
            .I(N__43550));
    CEMux I__9932 (
            .O(N__43572),
            .I(N__43550));
    CEMux I__9931 (
            .O(N__43571),
            .I(N__43550));
    CEMux I__9930 (
            .O(N__43570),
            .I(N__43550));
    CEMux I__9929 (
            .O(N__43569),
            .I(N__43550));
    CEMux I__9928 (
            .O(N__43568),
            .I(N__43550));
    CEMux I__9927 (
            .O(N__43567),
            .I(N__43550));
    GlobalMux I__9926 (
            .O(N__43550),
            .I(N__43547));
    gio2CtrlBuf I__9925 (
            .O(N__43547),
            .I(\current_shift_inst.timer_s1.N_162_i_g ));
    InMux I__9924 (
            .O(N__43544),
            .I(N__43541));
    LocalMux I__9923 (
            .O(N__43541),
            .I(N__43538));
    Span4Mux_h I__9922 (
            .O(N__43538),
            .I(N__43535));
    Odrv4 I__9921 (
            .O(N__43535),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    InMux I__9920 (
            .O(N__43532),
            .I(N__43529));
    LocalMux I__9919 (
            .O(N__43529),
            .I(N__43526));
    Span4Mux_h I__9918 (
            .O(N__43526),
            .I(N__43523));
    Odrv4 I__9917 (
            .O(N__43523),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    CascadeMux I__9916 (
            .O(N__43520),
            .I(N__43517));
    InMux I__9915 (
            .O(N__43517),
            .I(N__43513));
    InMux I__9914 (
            .O(N__43516),
            .I(N__43510));
    LocalMux I__9913 (
            .O(N__43513),
            .I(N__43507));
    LocalMux I__9912 (
            .O(N__43510),
            .I(N__43501));
    Span4Mux_h I__9911 (
            .O(N__43507),
            .I(N__43501));
    InMux I__9910 (
            .O(N__43506),
            .I(N__43498));
    Odrv4 I__9909 (
            .O(N__43501),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__9908 (
            .O(N__43498),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__9907 (
            .O(N__43493),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__9906 (
            .O(N__43490),
            .I(N__43487));
    LocalMux I__9905 (
            .O(N__43487),
            .I(N__43484));
    Span4Mux_v I__9904 (
            .O(N__43484),
            .I(N__43481));
    Odrv4 I__9903 (
            .O(N__43481),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__9902 (
            .O(N__43478),
            .I(N__43475));
    LocalMux I__9901 (
            .O(N__43475),
            .I(N__43470));
    InMux I__9900 (
            .O(N__43474),
            .I(N__43467));
    InMux I__9899 (
            .O(N__43473),
            .I(N__43464));
    Odrv4 I__9898 (
            .O(N__43470),
            .I(\current_shift_inst.un4_control_input1_22 ));
    LocalMux I__9897 (
            .O(N__43467),
            .I(\current_shift_inst.un4_control_input1_22 ));
    LocalMux I__9896 (
            .O(N__43464),
            .I(\current_shift_inst.un4_control_input1_22 ));
    InMux I__9895 (
            .O(N__43457),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__9894 (
            .O(N__43454),
            .I(N__43451));
    LocalMux I__9893 (
            .O(N__43451),
            .I(N__43448));
    Span4Mux_h I__9892 (
            .O(N__43448),
            .I(N__43445));
    Odrv4 I__9891 (
            .O(N__43445),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    CascadeMux I__9890 (
            .O(N__43442),
            .I(N__43438));
    InMux I__9889 (
            .O(N__43441),
            .I(N__43435));
    InMux I__9888 (
            .O(N__43438),
            .I(N__43432));
    LocalMux I__9887 (
            .O(N__43435),
            .I(N__43429));
    LocalMux I__9886 (
            .O(N__43432),
            .I(N__43424));
    Span4Mux_v I__9885 (
            .O(N__43429),
            .I(N__43424));
    Sp12to4 I__9884 (
            .O(N__43424),
            .I(N__43420));
    InMux I__9883 (
            .O(N__43423),
            .I(N__43417));
    Odrv12 I__9882 (
            .O(N__43420),
            .I(\current_shift_inst.un4_control_input1_23 ));
    LocalMux I__9881 (
            .O(N__43417),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__9880 (
            .O(N__43412),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__9879 (
            .O(N__43409),
            .I(N__43406));
    LocalMux I__9878 (
            .O(N__43406),
            .I(N__43403));
    Span4Mux_h I__9877 (
            .O(N__43403),
            .I(N__43400));
    Odrv4 I__9876 (
            .O(N__43400),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    CascadeMux I__9875 (
            .O(N__43397),
            .I(N__43393));
    InMux I__9874 (
            .O(N__43396),
            .I(N__43389));
    InMux I__9873 (
            .O(N__43393),
            .I(N__43386));
    InMux I__9872 (
            .O(N__43392),
            .I(N__43383));
    LocalMux I__9871 (
            .O(N__43389),
            .I(N__43378));
    LocalMux I__9870 (
            .O(N__43386),
            .I(N__43378));
    LocalMux I__9869 (
            .O(N__43383),
            .I(N__43375));
    Odrv12 I__9868 (
            .O(N__43378),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__9867 (
            .O(N__43375),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__9866 (
            .O(N__43370),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__9865 (
            .O(N__43367),
            .I(N__43364));
    LocalMux I__9864 (
            .O(N__43364),
            .I(N__43361));
    Span12Mux_v I__9863 (
            .O(N__43361),
            .I(N__43358));
    Odrv12 I__9862 (
            .O(N__43358),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    InMux I__9861 (
            .O(N__43355),
            .I(N__43352));
    LocalMux I__9860 (
            .O(N__43352),
            .I(N__43349));
    Span4Mux_h I__9859 (
            .O(N__43349),
            .I(N__43345));
    InMux I__9858 (
            .O(N__43348),
            .I(N__43342));
    Span4Mux_h I__9857 (
            .O(N__43345),
            .I(N__43338));
    LocalMux I__9856 (
            .O(N__43342),
            .I(N__43335));
    InMux I__9855 (
            .O(N__43341),
            .I(N__43332));
    Odrv4 I__9854 (
            .O(N__43338),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv4 I__9853 (
            .O(N__43335),
            .I(\current_shift_inst.un4_control_input1_25 ));
    LocalMux I__9852 (
            .O(N__43332),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__9851 (
            .O(N__43325),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__9850 (
            .O(N__43322),
            .I(N__43319));
    LocalMux I__9849 (
            .O(N__43319),
            .I(N__43316));
    Span4Mux_h I__9848 (
            .O(N__43316),
            .I(N__43313));
    Odrv4 I__9847 (
            .O(N__43313),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    CascadeMux I__9846 (
            .O(N__43310),
            .I(N__43306));
    CascadeMux I__9845 (
            .O(N__43309),
            .I(N__43303));
    InMux I__9844 (
            .O(N__43306),
            .I(N__43300));
    InMux I__9843 (
            .O(N__43303),
            .I(N__43297));
    LocalMux I__9842 (
            .O(N__43300),
            .I(N__43294));
    LocalMux I__9841 (
            .O(N__43297),
            .I(N__43291));
    Sp12to4 I__9840 (
            .O(N__43294),
            .I(N__43285));
    Span12Mux_h I__9839 (
            .O(N__43291),
            .I(N__43285));
    InMux I__9838 (
            .O(N__43290),
            .I(N__43282));
    Odrv12 I__9837 (
            .O(N__43285),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__9836 (
            .O(N__43282),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__9835 (
            .O(N__43277),
            .I(bfn_18_17_0_));
    InMux I__9834 (
            .O(N__43274),
            .I(N__43271));
    LocalMux I__9833 (
            .O(N__43271),
            .I(N__43268));
    Span4Mux_h I__9832 (
            .O(N__43268),
            .I(N__43265));
    Odrv4 I__9831 (
            .O(N__43265),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__9830 (
            .O(N__43262),
            .I(N__43258));
    InMux I__9829 (
            .O(N__43261),
            .I(N__43255));
    LocalMux I__9828 (
            .O(N__43258),
            .I(N__43252));
    LocalMux I__9827 (
            .O(N__43255),
            .I(N__43249));
    Span4Mux_h I__9826 (
            .O(N__43252),
            .I(N__43245));
    Span4Mux_v I__9825 (
            .O(N__43249),
            .I(N__43242));
    InMux I__9824 (
            .O(N__43248),
            .I(N__43239));
    Odrv4 I__9823 (
            .O(N__43245),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__9822 (
            .O(N__43242),
            .I(\current_shift_inst.un4_control_input1_27 ));
    LocalMux I__9821 (
            .O(N__43239),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__9820 (
            .O(N__43232),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__9819 (
            .O(N__43229),
            .I(N__43226));
    LocalMux I__9818 (
            .O(N__43226),
            .I(N__43223));
    Span4Mux_h I__9817 (
            .O(N__43223),
            .I(N__43220));
    Odrv4 I__9816 (
            .O(N__43220),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__9815 (
            .O(N__43217),
            .I(N__43211));
    InMux I__9814 (
            .O(N__43216),
            .I(N__43211));
    LocalMux I__9813 (
            .O(N__43211),
            .I(N__43207));
    InMux I__9812 (
            .O(N__43210),
            .I(N__43204));
    Odrv4 I__9811 (
            .O(N__43207),
            .I(\current_shift_inst.un4_control_input1_28 ));
    LocalMux I__9810 (
            .O(N__43204),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__9809 (
            .O(N__43199),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__9808 (
            .O(N__43196),
            .I(N__43193));
    LocalMux I__9807 (
            .O(N__43193),
            .I(N__43190));
    Span4Mux_h I__9806 (
            .O(N__43190),
            .I(N__43187));
    Odrv4 I__9805 (
            .O(N__43187),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__9804 (
            .O(N__43184),
            .I(N__43178));
    InMux I__9803 (
            .O(N__43183),
            .I(N__43178));
    LocalMux I__9802 (
            .O(N__43178),
            .I(N__43174));
    InMux I__9801 (
            .O(N__43177),
            .I(N__43171));
    Odrv12 I__9800 (
            .O(N__43174),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__9799 (
            .O(N__43171),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__9798 (
            .O(N__43166),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__9797 (
            .O(N__43163),
            .I(N__43160));
    LocalMux I__9796 (
            .O(N__43160),
            .I(N__43157));
    Span12Mux_v I__9795 (
            .O(N__43157),
            .I(N__43154));
    Odrv12 I__9794 (
            .O(N__43154),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__9793 (
            .O(N__43151),
            .I(N__43148));
    LocalMux I__9792 (
            .O(N__43148),
            .I(N__43144));
    InMux I__9791 (
            .O(N__43147),
            .I(N__43141));
    Span4Mux_h I__9790 (
            .O(N__43144),
            .I(N__43137));
    LocalMux I__9789 (
            .O(N__43141),
            .I(N__43134));
    InMux I__9788 (
            .O(N__43140),
            .I(N__43131));
    Odrv4 I__9787 (
            .O(N__43137),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv12 I__9786 (
            .O(N__43134),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__9785 (
            .O(N__43131),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__9784 (
            .O(N__43124),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    CascadeMux I__9783 (
            .O(N__43121),
            .I(N__43118));
    InMux I__9782 (
            .O(N__43118),
            .I(N__43114));
    CascadeMux I__9781 (
            .O(N__43117),
            .I(N__43111));
    LocalMux I__9780 (
            .O(N__43114),
            .I(N__43108));
    InMux I__9779 (
            .O(N__43111),
            .I(N__43105));
    Span4Mux_v I__9778 (
            .O(N__43108),
            .I(N__43102));
    LocalMux I__9777 (
            .O(N__43105),
            .I(N__43098));
    Span4Mux_h I__9776 (
            .O(N__43102),
            .I(N__43095));
    InMux I__9775 (
            .O(N__43101),
            .I(N__43092));
    Odrv4 I__9774 (
            .O(N__43098),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__9773 (
            .O(N__43095),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__9772 (
            .O(N__43092),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__9771 (
            .O(N__43085),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__9770 (
            .O(N__43082),
            .I(N__43079));
    LocalMux I__9769 (
            .O(N__43079),
            .I(N__43076));
    Span4Mux_h I__9768 (
            .O(N__43076),
            .I(N__43073));
    Odrv4 I__9767 (
            .O(N__43073),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__9766 (
            .O(N__43070),
            .I(N__43066));
    InMux I__9765 (
            .O(N__43069),
            .I(N__43063));
    LocalMux I__9764 (
            .O(N__43066),
            .I(N__43059));
    LocalMux I__9763 (
            .O(N__43063),
            .I(N__43056));
    InMux I__9762 (
            .O(N__43062),
            .I(N__43053));
    Odrv12 I__9761 (
            .O(N__43059),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__9760 (
            .O(N__43056),
            .I(\current_shift_inst.un4_control_input1_16 ));
    LocalMux I__9759 (
            .O(N__43053),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__9758 (
            .O(N__43046),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__9757 (
            .O(N__43043),
            .I(N__43040));
    LocalMux I__9756 (
            .O(N__43040),
            .I(N__43037));
    Span4Mux_h I__9755 (
            .O(N__43037),
            .I(N__43034));
    Odrv4 I__9754 (
            .O(N__43034),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__9753 (
            .O(N__43031),
            .I(N__43028));
    LocalMux I__9752 (
            .O(N__43028),
            .I(N__43024));
    InMux I__9751 (
            .O(N__43027),
            .I(N__43021));
    Span4Mux_h I__9750 (
            .O(N__43024),
            .I(N__43018));
    LocalMux I__9749 (
            .O(N__43021),
            .I(N__43014));
    Span4Mux_h I__9748 (
            .O(N__43018),
            .I(N__43011));
    InMux I__9747 (
            .O(N__43017),
            .I(N__43008));
    Odrv4 I__9746 (
            .O(N__43014),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__9745 (
            .O(N__43011),
            .I(\current_shift_inst.un4_control_input1_17 ));
    LocalMux I__9744 (
            .O(N__43008),
            .I(\current_shift_inst.un4_control_input1_17 ));
    InMux I__9743 (
            .O(N__43001),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__9742 (
            .O(N__42998),
            .I(N__42995));
    LocalMux I__9741 (
            .O(N__42995),
            .I(N__42990));
    CascadeMux I__9740 (
            .O(N__42994),
            .I(N__42987));
    InMux I__9739 (
            .O(N__42993),
            .I(N__42984));
    Span4Mux_h I__9738 (
            .O(N__42990),
            .I(N__42981));
    InMux I__9737 (
            .O(N__42987),
            .I(N__42978));
    LocalMux I__9736 (
            .O(N__42984),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__9735 (
            .O(N__42981),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__9734 (
            .O(N__42978),
            .I(\current_shift_inst.un4_control_input1_18 ));
    InMux I__9733 (
            .O(N__42971),
            .I(bfn_18_16_0_));
    InMux I__9732 (
            .O(N__42968),
            .I(N__42965));
    LocalMux I__9731 (
            .O(N__42965),
            .I(N__42962));
    Span4Mux_h I__9730 (
            .O(N__42962),
            .I(N__42959));
    Odrv4 I__9729 (
            .O(N__42959),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__9728 (
            .O(N__42956),
            .I(N__42952));
    InMux I__9727 (
            .O(N__42955),
            .I(N__42949));
    LocalMux I__9726 (
            .O(N__42952),
            .I(N__42943));
    LocalMux I__9725 (
            .O(N__42949),
            .I(N__42943));
    InMux I__9724 (
            .O(N__42948),
            .I(N__42940));
    Odrv12 I__9723 (
            .O(N__42943),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__9722 (
            .O(N__42940),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__9721 (
            .O(N__42935),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    CascadeMux I__9720 (
            .O(N__42932),
            .I(N__42928));
    InMux I__9719 (
            .O(N__42931),
            .I(N__42924));
    InMux I__9718 (
            .O(N__42928),
            .I(N__42921));
    InMux I__9717 (
            .O(N__42927),
            .I(N__42918));
    LocalMux I__9716 (
            .O(N__42924),
            .I(N__42915));
    LocalMux I__9715 (
            .O(N__42921),
            .I(N__42910));
    LocalMux I__9714 (
            .O(N__42918),
            .I(N__42910));
    Odrv12 I__9713 (
            .O(N__42915),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__9712 (
            .O(N__42910),
            .I(\current_shift_inst.un4_control_input1_20 ));
    InMux I__9711 (
            .O(N__42905),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__9710 (
            .O(N__42902),
            .I(N__42899));
    LocalMux I__9709 (
            .O(N__42899),
            .I(N__42896));
    Span4Mux_h I__9708 (
            .O(N__42896),
            .I(N__42893));
    Odrv4 I__9707 (
            .O(N__42893),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    CascadeMux I__9706 (
            .O(N__42890),
            .I(N__42886));
    CascadeMux I__9705 (
            .O(N__42889),
            .I(N__42883));
    InMux I__9704 (
            .O(N__42886),
            .I(N__42880));
    InMux I__9703 (
            .O(N__42883),
            .I(N__42877));
    LocalMux I__9702 (
            .O(N__42880),
            .I(N__42871));
    LocalMux I__9701 (
            .O(N__42877),
            .I(N__42871));
    InMux I__9700 (
            .O(N__42876),
            .I(N__42868));
    Odrv12 I__9699 (
            .O(N__42871),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__9698 (
            .O(N__42868),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__9697 (
            .O(N__42863),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__9696 (
            .O(N__42860),
            .I(N__42857));
    LocalMux I__9695 (
            .O(N__42857),
            .I(N__42854));
    Span4Mux_h I__9694 (
            .O(N__42854),
            .I(N__42851));
    Span4Mux_v I__9693 (
            .O(N__42851),
            .I(N__42848));
    Odrv4 I__9692 (
            .O(N__42848),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__9691 (
            .O(N__42845),
            .I(N__42839));
    InMux I__9690 (
            .O(N__42844),
            .I(N__42839));
    LocalMux I__9689 (
            .O(N__42839),
            .I(N__42835));
    InMux I__9688 (
            .O(N__42838),
            .I(N__42832));
    Odrv4 I__9687 (
            .O(N__42835),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__9686 (
            .O(N__42832),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__9685 (
            .O(N__42827),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__9684 (
            .O(N__42824),
            .I(N__42821));
    LocalMux I__9683 (
            .O(N__42821),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__9682 (
            .O(N__42818),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__9681 (
            .O(N__42815),
            .I(N__42812));
    LocalMux I__9680 (
            .O(N__42812),
            .I(N__42809));
    Span12Mux_v I__9679 (
            .O(N__42809),
            .I(N__42806));
    Odrv12 I__9678 (
            .O(N__42806),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__9677 (
            .O(N__42803),
            .I(N__42800));
    LocalMux I__9676 (
            .O(N__42800),
            .I(N__42796));
    InMux I__9675 (
            .O(N__42799),
            .I(N__42793));
    Span4Mux_h I__9674 (
            .O(N__42796),
            .I(N__42789));
    LocalMux I__9673 (
            .O(N__42793),
            .I(N__42786));
    InMux I__9672 (
            .O(N__42792),
            .I(N__42783));
    Odrv4 I__9671 (
            .O(N__42789),
            .I(\current_shift_inst.un4_control_input1_8 ));
    Odrv12 I__9670 (
            .O(N__42786),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__9669 (
            .O(N__42783),
            .I(\current_shift_inst.un4_control_input1_8 ));
    InMux I__9668 (
            .O(N__42776),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__9667 (
            .O(N__42773),
            .I(N__42770));
    LocalMux I__9666 (
            .O(N__42770),
            .I(N__42767));
    Span4Mux_v I__9665 (
            .O(N__42767),
            .I(N__42764));
    Odrv4 I__9664 (
            .O(N__42764),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__9663 (
            .O(N__42761),
            .I(N__42757));
    CascadeMux I__9662 (
            .O(N__42760),
            .I(N__42754));
    LocalMux I__9661 (
            .O(N__42757),
            .I(N__42751));
    InMux I__9660 (
            .O(N__42754),
            .I(N__42748));
    Span4Mux_v I__9659 (
            .O(N__42751),
            .I(N__42742));
    LocalMux I__9658 (
            .O(N__42748),
            .I(N__42742));
    InMux I__9657 (
            .O(N__42747),
            .I(N__42739));
    Odrv4 I__9656 (
            .O(N__42742),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__9655 (
            .O(N__42739),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__9654 (
            .O(N__42734),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__9653 (
            .O(N__42731),
            .I(N__42728));
    LocalMux I__9652 (
            .O(N__42728),
            .I(N__42725));
    Span4Mux_h I__9651 (
            .O(N__42725),
            .I(N__42722));
    Odrv4 I__9650 (
            .O(N__42722),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    CascadeMux I__9649 (
            .O(N__42719),
            .I(N__42716));
    InMux I__9648 (
            .O(N__42716),
            .I(N__42712));
    InMux I__9647 (
            .O(N__42715),
            .I(N__42709));
    LocalMux I__9646 (
            .O(N__42712),
            .I(N__42706));
    LocalMux I__9645 (
            .O(N__42709),
            .I(N__42703));
    Span4Mux_h I__9644 (
            .O(N__42706),
            .I(N__42697));
    Span4Mux_h I__9643 (
            .O(N__42703),
            .I(N__42697));
    InMux I__9642 (
            .O(N__42702),
            .I(N__42694));
    Odrv4 I__9641 (
            .O(N__42697),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__9640 (
            .O(N__42694),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__9639 (
            .O(N__42689),
            .I(bfn_18_15_0_));
    InMux I__9638 (
            .O(N__42686),
            .I(N__42683));
    LocalMux I__9637 (
            .O(N__42683),
            .I(N__42680));
    Span4Mux_h I__9636 (
            .O(N__42680),
            .I(N__42677));
    Span4Mux_h I__9635 (
            .O(N__42677),
            .I(N__42674));
    Odrv4 I__9634 (
            .O(N__42674),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    CascadeMux I__9633 (
            .O(N__42671),
            .I(N__42667));
    InMux I__9632 (
            .O(N__42670),
            .I(N__42664));
    InMux I__9631 (
            .O(N__42667),
            .I(N__42661));
    LocalMux I__9630 (
            .O(N__42664),
            .I(N__42655));
    LocalMux I__9629 (
            .O(N__42661),
            .I(N__42655));
    InMux I__9628 (
            .O(N__42660),
            .I(N__42652));
    Odrv12 I__9627 (
            .O(N__42655),
            .I(\current_shift_inst.un4_control_input1_11 ));
    LocalMux I__9626 (
            .O(N__42652),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__9625 (
            .O(N__42647),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__9624 (
            .O(N__42644),
            .I(N__42641));
    LocalMux I__9623 (
            .O(N__42641),
            .I(N__42638));
    Span4Mux_v I__9622 (
            .O(N__42638),
            .I(N__42635));
    Odrv4 I__9621 (
            .O(N__42635),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__9620 (
            .O(N__42632),
            .I(N__42628));
    InMux I__9619 (
            .O(N__42631),
            .I(N__42625));
    LocalMux I__9618 (
            .O(N__42628),
            .I(N__42622));
    LocalMux I__9617 (
            .O(N__42625),
            .I(N__42618));
    Span4Mux_h I__9616 (
            .O(N__42622),
            .I(N__42615));
    InMux I__9615 (
            .O(N__42621),
            .I(N__42612));
    Odrv12 I__9614 (
            .O(N__42618),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__9613 (
            .O(N__42615),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__9612 (
            .O(N__42612),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__9611 (
            .O(N__42605),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    CascadeMux I__9610 (
            .O(N__42602),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_));
    InMux I__9609 (
            .O(N__42599),
            .I(N__42593));
    InMux I__9608 (
            .O(N__42598),
            .I(N__42588));
    InMux I__9607 (
            .O(N__42597),
            .I(N__42588));
    InMux I__9606 (
            .O(N__42596),
            .I(N__42585));
    LocalMux I__9605 (
            .O(N__42593),
            .I(N__42582));
    LocalMux I__9604 (
            .O(N__42588),
            .I(N__42579));
    LocalMux I__9603 (
            .O(N__42585),
            .I(N__42576));
    Span4Mux_v I__9602 (
            .O(N__42582),
            .I(N__42573));
    Span4Mux_h I__9601 (
            .O(N__42579),
            .I(N__42570));
    Span12Mux_s10_h I__9600 (
            .O(N__42576),
            .I(N__42567));
    Odrv4 I__9599 (
            .O(N__42573),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv4 I__9598 (
            .O(N__42570),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv12 I__9597 (
            .O(N__42567),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__9596 (
            .O(N__42560),
            .I(N__42554));
    InMux I__9595 (
            .O(N__42559),
            .I(N__42554));
    LocalMux I__9594 (
            .O(N__42554),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    InMux I__9593 (
            .O(N__42551),
            .I(N__42548));
    LocalMux I__9592 (
            .O(N__42548),
            .I(N__42542));
    InMux I__9591 (
            .O(N__42547),
            .I(N__42537));
    InMux I__9590 (
            .O(N__42546),
            .I(N__42537));
    InMux I__9589 (
            .O(N__42545),
            .I(N__42534));
    Span4Mux_v I__9588 (
            .O(N__42542),
            .I(N__42529));
    LocalMux I__9587 (
            .O(N__42537),
            .I(N__42529));
    LocalMux I__9586 (
            .O(N__42534),
            .I(N__42526));
    Span4Mux_h I__9585 (
            .O(N__42529),
            .I(N__42523));
    Odrv12 I__9584 (
            .O(N__42526),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    Odrv4 I__9583 (
            .O(N__42523),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__9582 (
            .O(N__42518),
            .I(N__42514));
    InMux I__9581 (
            .O(N__42517),
            .I(N__42511));
    LocalMux I__9580 (
            .O(N__42514),
            .I(N__42507));
    LocalMux I__9579 (
            .O(N__42511),
            .I(N__42504));
    InMux I__9578 (
            .O(N__42510),
            .I(N__42501));
    Span4Mux_h I__9577 (
            .O(N__42507),
            .I(N__42498));
    Span4Mux_v I__9576 (
            .O(N__42504),
            .I(N__42495));
    LocalMux I__9575 (
            .O(N__42501),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv4 I__9574 (
            .O(N__42498),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv4 I__9573 (
            .O(N__42495),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    InMux I__9572 (
            .O(N__42488),
            .I(N__42485));
    LocalMux I__9571 (
            .O(N__42485),
            .I(N__42482));
    Odrv4 I__9570 (
            .O(N__42482),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__9569 (
            .O(N__42479),
            .I(N__42476));
    LocalMux I__9568 (
            .O(N__42476),
            .I(N__42473));
    Span4Mux_v I__9567 (
            .O(N__42473),
            .I(N__42470));
    Odrv4 I__9566 (
            .O(N__42470),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__9565 (
            .O(N__42467),
            .I(N__42463));
    InMux I__9564 (
            .O(N__42466),
            .I(N__42459));
    LocalMux I__9563 (
            .O(N__42463),
            .I(N__42456));
    InMux I__9562 (
            .O(N__42462),
            .I(N__42453));
    LocalMux I__9561 (
            .O(N__42459),
            .I(N__42450));
    Span4Mux_v I__9560 (
            .O(N__42456),
            .I(N__42445));
    LocalMux I__9559 (
            .O(N__42453),
            .I(N__42445));
    Span4Mux_h I__9558 (
            .O(N__42450),
            .I(N__42441));
    Span4Mux_h I__9557 (
            .O(N__42445),
            .I(N__42438));
    InMux I__9556 (
            .O(N__42444),
            .I(N__42435));
    Odrv4 I__9555 (
            .O(N__42441),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__9554 (
            .O(N__42438),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__9553 (
            .O(N__42435),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__9552 (
            .O(N__42428),
            .I(N__42425));
    LocalMux I__9551 (
            .O(N__42425),
            .I(N__42422));
    Span4Mux_h I__9550 (
            .O(N__42422),
            .I(N__42419));
    Odrv4 I__9549 (
            .O(N__42419),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__9548 (
            .O(N__42416),
            .I(N__42411));
    InMux I__9547 (
            .O(N__42415),
            .I(N__42408));
    InMux I__9546 (
            .O(N__42414),
            .I(N__42405));
    LocalMux I__9545 (
            .O(N__42411),
            .I(N__42400));
    LocalMux I__9544 (
            .O(N__42408),
            .I(N__42400));
    LocalMux I__9543 (
            .O(N__42405),
            .I(N__42397));
    Span4Mux_v I__9542 (
            .O(N__42400),
            .I(N__42394));
    Span12Mux_s10_h I__9541 (
            .O(N__42397),
            .I(N__42391));
    Span4Mux_v I__9540 (
            .O(N__42394),
            .I(N__42388));
    Odrv12 I__9539 (
            .O(N__42391),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__9538 (
            .O(N__42388),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    InMux I__9537 (
            .O(N__42383),
            .I(N__42377));
    InMux I__9536 (
            .O(N__42382),
            .I(N__42374));
    InMux I__9535 (
            .O(N__42381),
            .I(N__42371));
    InMux I__9534 (
            .O(N__42380),
            .I(N__42355));
    LocalMux I__9533 (
            .O(N__42377),
            .I(N__42352));
    LocalMux I__9532 (
            .O(N__42374),
            .I(N__42349));
    LocalMux I__9531 (
            .O(N__42371),
            .I(N__42346));
    InMux I__9530 (
            .O(N__42370),
            .I(N__42331));
    InMux I__9529 (
            .O(N__42369),
            .I(N__42331));
    InMux I__9528 (
            .O(N__42368),
            .I(N__42331));
    InMux I__9527 (
            .O(N__42367),
            .I(N__42331));
    InMux I__9526 (
            .O(N__42366),
            .I(N__42331));
    InMux I__9525 (
            .O(N__42365),
            .I(N__42331));
    InMux I__9524 (
            .O(N__42364),
            .I(N__42331));
    InMux I__9523 (
            .O(N__42363),
            .I(N__42318));
    InMux I__9522 (
            .O(N__42362),
            .I(N__42318));
    InMux I__9521 (
            .O(N__42361),
            .I(N__42318));
    InMux I__9520 (
            .O(N__42360),
            .I(N__42318));
    InMux I__9519 (
            .O(N__42359),
            .I(N__42318));
    InMux I__9518 (
            .O(N__42358),
            .I(N__42318));
    LocalMux I__9517 (
            .O(N__42355),
            .I(N__42305));
    Span4Mux_h I__9516 (
            .O(N__42352),
            .I(N__42305));
    Span4Mux_v I__9515 (
            .O(N__42349),
            .I(N__42296));
    Span4Mux_h I__9514 (
            .O(N__42346),
            .I(N__42296));
    LocalMux I__9513 (
            .O(N__42331),
            .I(N__42296));
    LocalMux I__9512 (
            .O(N__42318),
            .I(N__42296));
    InMux I__9511 (
            .O(N__42317),
            .I(N__42287));
    InMux I__9510 (
            .O(N__42316),
            .I(N__42287));
    InMux I__9509 (
            .O(N__42315),
            .I(N__42287));
    InMux I__9508 (
            .O(N__42314),
            .I(N__42287));
    InMux I__9507 (
            .O(N__42313),
            .I(N__42278));
    InMux I__9506 (
            .O(N__42312),
            .I(N__42278));
    InMux I__9505 (
            .O(N__42311),
            .I(N__42278));
    InMux I__9504 (
            .O(N__42310),
            .I(N__42278));
    Span4Mux_h I__9503 (
            .O(N__42305),
            .I(N__42275));
    Odrv4 I__9502 (
            .O(N__42296),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__9501 (
            .O(N__42287),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__9500 (
            .O(N__42278),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__9499 (
            .O(N__42275),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    CascadeMux I__9498 (
            .O(N__42266),
            .I(N__42262));
    InMux I__9497 (
            .O(N__42265),
            .I(N__42258));
    InMux I__9496 (
            .O(N__42262),
            .I(N__42255));
    InMux I__9495 (
            .O(N__42261),
            .I(N__42252));
    LocalMux I__9494 (
            .O(N__42258),
            .I(N__42247));
    LocalMux I__9493 (
            .O(N__42255),
            .I(N__42247));
    LocalMux I__9492 (
            .O(N__42252),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    Odrv12 I__9491 (
            .O(N__42247),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__9490 (
            .O(N__42242),
            .I(N__42239));
    LocalMux I__9489 (
            .O(N__42239),
            .I(N__42236));
    Span4Mux_h I__9488 (
            .O(N__42236),
            .I(N__42233));
    Span4Mux_v I__9487 (
            .O(N__42233),
            .I(N__42230));
    Odrv4 I__9486 (
            .O(N__42230),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__9485 (
            .O(N__42227),
            .I(N__42221));
    InMux I__9484 (
            .O(N__42226),
            .I(N__42221));
    LocalMux I__9483 (
            .O(N__42221),
            .I(N__42218));
    Span4Mux_h I__9482 (
            .O(N__42218),
            .I(N__42214));
    InMux I__9481 (
            .O(N__42217),
            .I(N__42211));
    Odrv4 I__9480 (
            .O(N__42214),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__9479 (
            .O(N__42211),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__9478 (
            .O(N__42206),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__9477 (
            .O(N__42203),
            .I(N__42200));
    LocalMux I__9476 (
            .O(N__42200),
            .I(N__42197));
    Span4Mux_h I__9475 (
            .O(N__42197),
            .I(N__42194));
    Odrv4 I__9474 (
            .O(N__42194),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__9473 (
            .O(N__42191),
            .I(N__42187));
    InMux I__9472 (
            .O(N__42190),
            .I(N__42184));
    LocalMux I__9471 (
            .O(N__42187),
            .I(N__42181));
    LocalMux I__9470 (
            .O(N__42184),
            .I(N__42178));
    Span4Mux_v I__9469 (
            .O(N__42181),
            .I(N__42172));
    Span4Mux_h I__9468 (
            .O(N__42178),
            .I(N__42172));
    InMux I__9467 (
            .O(N__42177),
            .I(N__42169));
    Odrv4 I__9466 (
            .O(N__42172),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__9465 (
            .O(N__42169),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__9464 (
            .O(N__42164),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    CascadeMux I__9463 (
            .O(N__42161),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ));
    CascadeMux I__9462 (
            .O(N__42158),
            .I(N__42155));
    InMux I__9461 (
            .O(N__42155),
            .I(N__42152));
    LocalMux I__9460 (
            .O(N__42152),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ));
    CascadeMux I__9459 (
            .O(N__42149),
            .I(N__42146));
    InMux I__9458 (
            .O(N__42146),
            .I(N__42142));
    InMux I__9457 (
            .O(N__42145),
            .I(N__42139));
    LocalMux I__9456 (
            .O(N__42142),
            .I(N__42136));
    LocalMux I__9455 (
            .O(N__42139),
            .I(N__42133));
    Span4Mux_h I__9454 (
            .O(N__42136),
            .I(N__42130));
    Span12Mux_v I__9453 (
            .O(N__42133),
            .I(N__42127));
    Odrv4 I__9452 (
            .O(N__42130),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv12 I__9451 (
            .O(N__42127),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__9450 (
            .O(N__42122),
            .I(N__42118));
    InMux I__9449 (
            .O(N__42121),
            .I(N__42115));
    LocalMux I__9448 (
            .O(N__42118),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    LocalMux I__9447 (
            .O(N__42115),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    InMux I__9446 (
            .O(N__42110),
            .I(N__42106));
    InMux I__9445 (
            .O(N__42109),
            .I(N__42103));
    LocalMux I__9444 (
            .O(N__42106),
            .I(N__42100));
    LocalMux I__9443 (
            .O(N__42103),
            .I(N__42097));
    Span4Mux_h I__9442 (
            .O(N__42100),
            .I(N__42094));
    Span4Mux_v I__9441 (
            .O(N__42097),
            .I(N__42091));
    Odrv4 I__9440 (
            .O(N__42094),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    Odrv4 I__9439 (
            .O(N__42091),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    CascadeMux I__9438 (
            .O(N__42086),
            .I(N__42083));
    InMux I__9437 (
            .O(N__42083),
            .I(N__42080));
    LocalMux I__9436 (
            .O(N__42080),
            .I(N__42077));
    Odrv4 I__9435 (
            .O(N__42077),
            .I(\phase_controller_inst1.stoper_tr.un4_running_df30 ));
    InMux I__9434 (
            .O(N__42074),
            .I(N__42071));
    LocalMux I__9433 (
            .O(N__42071),
            .I(N__42068));
    Span4Mux_h I__9432 (
            .O(N__42068),
            .I(N__42065));
    Odrv4 I__9431 (
            .O(N__42065),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ));
    InMux I__9430 (
            .O(N__42062),
            .I(N__42059));
    LocalMux I__9429 (
            .O(N__42059),
            .I(N__42055));
    InMux I__9428 (
            .O(N__42058),
            .I(N__42052));
    Odrv12 I__9427 (
            .O(N__42055),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__9426 (
            .O(N__42052),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__9425 (
            .O(N__42047),
            .I(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__9424 (
            .O(N__42044),
            .I(N__42041));
    LocalMux I__9423 (
            .O(N__42041),
            .I(N__42037));
    InMux I__9422 (
            .O(N__42040),
            .I(N__42034));
    Span4Mux_v I__9421 (
            .O(N__42037),
            .I(N__42031));
    LocalMux I__9420 (
            .O(N__42034),
            .I(N__42028));
    Span4Mux_v I__9419 (
            .O(N__42031),
            .I(N__42025));
    Span4Mux_v I__9418 (
            .O(N__42028),
            .I(N__42022));
    Span4Mux_h I__9417 (
            .O(N__42025),
            .I(N__42017));
    Span4Mux_h I__9416 (
            .O(N__42022),
            .I(N__42014));
    InMux I__9415 (
            .O(N__42021),
            .I(N__42009));
    InMux I__9414 (
            .O(N__42020),
            .I(N__42009));
    Odrv4 I__9413 (
            .O(N__42017),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    Odrv4 I__9412 (
            .O(N__42014),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    LocalMux I__9411 (
            .O(N__42009),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__9410 (
            .O(N__42002),
            .I(N__41999));
    LocalMux I__9409 (
            .O(N__41999),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ));
    InMux I__9408 (
            .O(N__41996),
            .I(N__41993));
    LocalMux I__9407 (
            .O(N__41993),
            .I(N__41990));
    Span4Mux_h I__9406 (
            .O(N__41990),
            .I(N__41987));
    Odrv4 I__9405 (
            .O(N__41987),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__9404 (
            .O(N__41984),
            .I(N__41979));
    InMux I__9403 (
            .O(N__41983),
            .I(N__41974));
    InMux I__9402 (
            .O(N__41982),
            .I(N__41974));
    LocalMux I__9401 (
            .O(N__41979),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    LocalMux I__9400 (
            .O(N__41974),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__9399 (
            .O(N__41969),
            .I(N__41965));
    InMux I__9398 (
            .O(N__41968),
            .I(N__41961));
    InMux I__9397 (
            .O(N__41965),
            .I(N__41956));
    InMux I__9396 (
            .O(N__41964),
            .I(N__41956));
    LocalMux I__9395 (
            .O(N__41961),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    LocalMux I__9394 (
            .O(N__41956),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    CascadeMux I__9393 (
            .O(N__41951),
            .I(N__41948));
    InMux I__9392 (
            .O(N__41948),
            .I(N__41945));
    LocalMux I__9391 (
            .O(N__41945),
            .I(N__41942));
    Span4Mux_h I__9390 (
            .O(N__41942),
            .I(N__41939));
    Odrv4 I__9389 (
            .O(N__41939),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    InMux I__9388 (
            .O(N__41936),
            .I(N__41932));
    CascadeMux I__9387 (
            .O(N__41935),
            .I(N__41929));
    LocalMux I__9386 (
            .O(N__41932),
            .I(N__41926));
    InMux I__9385 (
            .O(N__41929),
            .I(N__41922));
    Span4Mux_v I__9384 (
            .O(N__41926),
            .I(N__41919));
    InMux I__9383 (
            .O(N__41925),
            .I(N__41916));
    LocalMux I__9382 (
            .O(N__41922),
            .I(N__41911));
    Span4Mux_h I__9381 (
            .O(N__41919),
            .I(N__41911));
    LocalMux I__9380 (
            .O(N__41916),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    Odrv4 I__9379 (
            .O(N__41911),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    InMux I__9378 (
            .O(N__41906),
            .I(N__41901));
    InMux I__9377 (
            .O(N__41905),
            .I(N__41897));
    InMux I__9376 (
            .O(N__41904),
            .I(N__41894));
    LocalMux I__9375 (
            .O(N__41901),
            .I(N__41891));
    InMux I__9374 (
            .O(N__41900),
            .I(N__41888));
    LocalMux I__9373 (
            .O(N__41897),
            .I(N__41885));
    LocalMux I__9372 (
            .O(N__41894),
            .I(N__41880));
    Span4Mux_h I__9371 (
            .O(N__41891),
            .I(N__41880));
    LocalMux I__9370 (
            .O(N__41888),
            .I(N__41877));
    Span4Mux_h I__9369 (
            .O(N__41885),
            .I(N__41872));
    Span4Mux_v I__9368 (
            .O(N__41880),
            .I(N__41872));
    Odrv4 I__9367 (
            .O(N__41877),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__9366 (
            .O(N__41872),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    CascadeMux I__9365 (
            .O(N__41867),
            .I(N__41864));
    InMux I__9364 (
            .O(N__41864),
            .I(N__41858));
    InMux I__9363 (
            .O(N__41863),
            .I(N__41858));
    LocalMux I__9362 (
            .O(N__41858),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__9361 (
            .O(N__41855),
            .I(N__41852));
    LocalMux I__9360 (
            .O(N__41852),
            .I(N__41849));
    Span4Mux_h I__9359 (
            .O(N__41849),
            .I(N__41846));
    Span4Mux_v I__9358 (
            .O(N__41846),
            .I(N__41842));
    InMux I__9357 (
            .O(N__41845),
            .I(N__41839));
    Odrv4 I__9356 (
            .O(N__41842),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    LocalMux I__9355 (
            .O(N__41839),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    InMux I__9354 (
            .O(N__41834),
            .I(N__41830));
    InMux I__9353 (
            .O(N__41833),
            .I(N__41826));
    LocalMux I__9352 (
            .O(N__41830),
            .I(N__41823));
    InMux I__9351 (
            .O(N__41829),
            .I(N__41820));
    LocalMux I__9350 (
            .O(N__41826),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    Odrv4 I__9349 (
            .O(N__41823),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    LocalMux I__9348 (
            .O(N__41820),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    InMux I__9347 (
            .O(N__41813),
            .I(N__41810));
    LocalMux I__9346 (
            .O(N__41810),
            .I(N__41805));
    InMux I__9345 (
            .O(N__41809),
            .I(N__41802));
    InMux I__9344 (
            .O(N__41808),
            .I(N__41799));
    Span4Mux_v I__9343 (
            .O(N__41805),
            .I(N__41792));
    LocalMux I__9342 (
            .O(N__41802),
            .I(N__41792));
    LocalMux I__9341 (
            .O(N__41799),
            .I(N__41792));
    Span4Mux_h I__9340 (
            .O(N__41792),
            .I(N__41788));
    InMux I__9339 (
            .O(N__41791),
            .I(N__41785));
    Odrv4 I__9338 (
            .O(N__41788),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    LocalMux I__9337 (
            .O(N__41785),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    CascadeMux I__9336 (
            .O(N__41780),
            .I(N__41777));
    InMux I__9335 (
            .O(N__41777),
            .I(N__41774));
    LocalMux I__9334 (
            .O(N__41774),
            .I(N__41771));
    Span4Mux_v I__9333 (
            .O(N__41771),
            .I(N__41768));
    Odrv4 I__9332 (
            .O(N__41768),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    InMux I__9331 (
            .O(N__41765),
            .I(N__41761));
    InMux I__9330 (
            .O(N__41764),
            .I(N__41758));
    LocalMux I__9329 (
            .O(N__41761),
            .I(N__41755));
    LocalMux I__9328 (
            .O(N__41758),
            .I(N__41749));
    Span4Mux_v I__9327 (
            .O(N__41755),
            .I(N__41749));
    InMux I__9326 (
            .O(N__41754),
            .I(N__41746));
    Odrv4 I__9325 (
            .O(N__41749),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    LocalMux I__9324 (
            .O(N__41746),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    CascadeMux I__9323 (
            .O(N__41741),
            .I(N__41735));
    CascadeMux I__9322 (
            .O(N__41740),
            .I(N__41732));
    InMux I__9321 (
            .O(N__41739),
            .I(N__41729));
    InMux I__9320 (
            .O(N__41738),
            .I(N__41726));
    InMux I__9319 (
            .O(N__41735),
            .I(N__41723));
    InMux I__9318 (
            .O(N__41732),
            .I(N__41720));
    LocalMux I__9317 (
            .O(N__41729),
            .I(N__41717));
    LocalMux I__9316 (
            .O(N__41726),
            .I(N__41712));
    LocalMux I__9315 (
            .O(N__41723),
            .I(N__41712));
    LocalMux I__9314 (
            .O(N__41720),
            .I(N__41707));
    Span4Mux_h I__9313 (
            .O(N__41717),
            .I(N__41707));
    Span4Mux_h I__9312 (
            .O(N__41712),
            .I(N__41704));
    Span4Mux_v I__9311 (
            .O(N__41707),
            .I(N__41701));
    Span4Mux_v I__9310 (
            .O(N__41704),
            .I(N__41698));
    Odrv4 I__9309 (
            .O(N__41701),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv4 I__9308 (
            .O(N__41698),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__9307 (
            .O(N__41693),
            .I(N__41688));
    InMux I__9306 (
            .O(N__41692),
            .I(N__41685));
    InMux I__9305 (
            .O(N__41691),
            .I(N__41682));
    LocalMux I__9304 (
            .O(N__41688),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__9303 (
            .O(N__41685),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__9302 (
            .O(N__41682),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    InMux I__9301 (
            .O(N__41675),
            .I(N__41669));
    InMux I__9300 (
            .O(N__41674),
            .I(N__41666));
    InMux I__9299 (
            .O(N__41673),
            .I(N__41663));
    InMux I__9298 (
            .O(N__41672),
            .I(N__41660));
    LocalMux I__9297 (
            .O(N__41669),
            .I(N__41657));
    LocalMux I__9296 (
            .O(N__41666),
            .I(N__41652));
    LocalMux I__9295 (
            .O(N__41663),
            .I(N__41652));
    LocalMux I__9294 (
            .O(N__41660),
            .I(N__41649));
    Span4Mux_h I__9293 (
            .O(N__41657),
            .I(N__41644));
    Span4Mux_v I__9292 (
            .O(N__41652),
            .I(N__41644));
    Span4Mux_h I__9291 (
            .O(N__41649),
            .I(N__41641));
    Span4Mux_v I__9290 (
            .O(N__41644),
            .I(N__41638));
    Span4Mux_v I__9289 (
            .O(N__41641),
            .I(N__41635));
    Odrv4 I__9288 (
            .O(N__41638),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    Odrv4 I__9287 (
            .O(N__41635),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__9286 (
            .O(N__41630),
            .I(N__41626));
    InMux I__9285 (
            .O(N__41629),
            .I(N__41623));
    LocalMux I__9284 (
            .O(N__41626),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    LocalMux I__9283 (
            .O(N__41623),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    CascadeMux I__9282 (
            .O(N__41618),
            .I(N__41615));
    InMux I__9281 (
            .O(N__41615),
            .I(N__41612));
    LocalMux I__9280 (
            .O(N__41612),
            .I(N__41609));
    Span4Mux_v I__9279 (
            .O(N__41609),
            .I(N__41606));
    Odrv4 I__9278 (
            .O(N__41606),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    InMux I__9277 (
            .O(N__41603),
            .I(N__41597));
    InMux I__9276 (
            .O(N__41602),
            .I(N__41597));
    LocalMux I__9275 (
            .O(N__41597),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__9274 (
            .O(N__41594),
            .I(N__41588));
    InMux I__9273 (
            .O(N__41593),
            .I(N__41588));
    LocalMux I__9272 (
            .O(N__41588),
            .I(N__41584));
    InMux I__9271 (
            .O(N__41587),
            .I(N__41581));
    Span4Mux_v I__9270 (
            .O(N__41584),
            .I(N__41578));
    LocalMux I__9269 (
            .O(N__41581),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__9268 (
            .O(N__41578),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    CascadeMux I__9267 (
            .O(N__41573),
            .I(N__41569));
    InMux I__9266 (
            .O(N__41572),
            .I(N__41563));
    InMux I__9265 (
            .O(N__41569),
            .I(N__41563));
    InMux I__9264 (
            .O(N__41568),
            .I(N__41560));
    LocalMux I__9263 (
            .O(N__41563),
            .I(N__41557));
    LocalMux I__9262 (
            .O(N__41560),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__9261 (
            .O(N__41557),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__9260 (
            .O(N__41552),
            .I(N__41548));
    InMux I__9259 (
            .O(N__41551),
            .I(N__41543));
    InMux I__9258 (
            .O(N__41548),
            .I(N__41543));
    LocalMux I__9257 (
            .O(N__41543),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__9256 (
            .O(N__41540),
            .I(N__41537));
    LocalMux I__9255 (
            .O(N__41537),
            .I(N__41534));
    Span4Mux_v I__9254 (
            .O(N__41534),
            .I(N__41531));
    Odrv4 I__9253 (
            .O(N__41531),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    InMux I__9252 (
            .O(N__41528),
            .I(N__41525));
    LocalMux I__9251 (
            .O(N__41525),
            .I(N__41521));
    InMux I__9250 (
            .O(N__41524),
            .I(N__41517));
    Span12Mux_h I__9249 (
            .O(N__41521),
            .I(N__41514));
    InMux I__9248 (
            .O(N__41520),
            .I(N__41511));
    LocalMux I__9247 (
            .O(N__41517),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    Odrv12 I__9246 (
            .O(N__41514),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    LocalMux I__9245 (
            .O(N__41511),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    InMux I__9244 (
            .O(N__41504),
            .I(N__41498));
    InMux I__9243 (
            .O(N__41503),
            .I(N__41495));
    InMux I__9242 (
            .O(N__41502),
            .I(N__41492));
    InMux I__9241 (
            .O(N__41501),
            .I(N__41489));
    LocalMux I__9240 (
            .O(N__41498),
            .I(N__41484));
    LocalMux I__9239 (
            .O(N__41495),
            .I(N__41484));
    LocalMux I__9238 (
            .O(N__41492),
            .I(N__41479));
    LocalMux I__9237 (
            .O(N__41489),
            .I(N__41479));
    Span4Mux_v I__9236 (
            .O(N__41484),
            .I(N__41474));
    Span4Mux_v I__9235 (
            .O(N__41479),
            .I(N__41474));
    Odrv4 I__9234 (
            .O(N__41474),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__9233 (
            .O(N__41471),
            .I(N__41468));
    LocalMux I__9232 (
            .O(N__41468),
            .I(N__41465));
    Span4Mux_h I__9231 (
            .O(N__41465),
            .I(N__41462));
    Odrv4 I__9230 (
            .O(N__41462),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    InMux I__9229 (
            .O(N__41459),
            .I(N__41456));
    LocalMux I__9228 (
            .O(N__41456),
            .I(N__41451));
    InMux I__9227 (
            .O(N__41455),
            .I(N__41448));
    InMux I__9226 (
            .O(N__41454),
            .I(N__41444));
    Span4Mux_v I__9225 (
            .O(N__41451),
            .I(N__41439));
    LocalMux I__9224 (
            .O(N__41448),
            .I(N__41439));
    InMux I__9223 (
            .O(N__41447),
            .I(N__41436));
    LocalMux I__9222 (
            .O(N__41444),
            .I(N__41433));
    Span4Mux_v I__9221 (
            .O(N__41439),
            .I(N__41428));
    LocalMux I__9220 (
            .O(N__41436),
            .I(N__41428));
    Span4Mux_v I__9219 (
            .O(N__41433),
            .I(N__41423));
    Span4Mux_h I__9218 (
            .O(N__41428),
            .I(N__41423));
    Odrv4 I__9217 (
            .O(N__41423),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__9216 (
            .O(N__41420),
            .I(N__41417));
    LocalMux I__9215 (
            .O(N__41417),
            .I(N__41412));
    InMux I__9214 (
            .O(N__41416),
            .I(N__41409));
    InMux I__9213 (
            .O(N__41415),
            .I(N__41406));
    Span4Mux_h I__9212 (
            .O(N__41412),
            .I(N__41401));
    LocalMux I__9211 (
            .O(N__41409),
            .I(N__41401));
    LocalMux I__9210 (
            .O(N__41406),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    Odrv4 I__9209 (
            .O(N__41401),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    InMux I__9208 (
            .O(N__41396),
            .I(N__41389));
    InMux I__9207 (
            .O(N__41395),
            .I(N__41389));
    InMux I__9206 (
            .O(N__41394),
            .I(N__41386));
    LocalMux I__9205 (
            .O(N__41389),
            .I(N__41383));
    LocalMux I__9204 (
            .O(N__41386),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__9203 (
            .O(N__41383),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__9202 (
            .O(N__41378),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    CascadeMux I__9201 (
            .O(N__41375),
            .I(N__41372));
    InMux I__9200 (
            .O(N__41372),
            .I(N__41368));
    InMux I__9199 (
            .O(N__41371),
            .I(N__41365));
    LocalMux I__9198 (
            .O(N__41368),
            .I(N__41362));
    LocalMux I__9197 (
            .O(N__41365),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__9196 (
            .O(N__41362),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__9195 (
            .O(N__41357),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__9194 (
            .O(N__41354),
            .I(N__41316));
    InMux I__9193 (
            .O(N__41353),
            .I(N__41316));
    InMux I__9192 (
            .O(N__41352),
            .I(N__41316));
    InMux I__9191 (
            .O(N__41351),
            .I(N__41316));
    InMux I__9190 (
            .O(N__41350),
            .I(N__41307));
    InMux I__9189 (
            .O(N__41349),
            .I(N__41307));
    InMux I__9188 (
            .O(N__41348),
            .I(N__41307));
    InMux I__9187 (
            .O(N__41347),
            .I(N__41307));
    InMux I__9186 (
            .O(N__41346),
            .I(N__41302));
    InMux I__9185 (
            .O(N__41345),
            .I(N__41302));
    InMux I__9184 (
            .O(N__41344),
            .I(N__41293));
    InMux I__9183 (
            .O(N__41343),
            .I(N__41293));
    InMux I__9182 (
            .O(N__41342),
            .I(N__41293));
    InMux I__9181 (
            .O(N__41341),
            .I(N__41293));
    InMux I__9180 (
            .O(N__41340),
            .I(N__41284));
    InMux I__9179 (
            .O(N__41339),
            .I(N__41284));
    InMux I__9178 (
            .O(N__41338),
            .I(N__41284));
    InMux I__9177 (
            .O(N__41337),
            .I(N__41284));
    InMux I__9176 (
            .O(N__41336),
            .I(N__41275));
    InMux I__9175 (
            .O(N__41335),
            .I(N__41275));
    InMux I__9174 (
            .O(N__41334),
            .I(N__41275));
    InMux I__9173 (
            .O(N__41333),
            .I(N__41275));
    InMux I__9172 (
            .O(N__41332),
            .I(N__41266));
    InMux I__9171 (
            .O(N__41331),
            .I(N__41266));
    InMux I__9170 (
            .O(N__41330),
            .I(N__41266));
    InMux I__9169 (
            .O(N__41329),
            .I(N__41266));
    InMux I__9168 (
            .O(N__41328),
            .I(N__41257));
    InMux I__9167 (
            .O(N__41327),
            .I(N__41257));
    InMux I__9166 (
            .O(N__41326),
            .I(N__41257));
    InMux I__9165 (
            .O(N__41325),
            .I(N__41257));
    LocalMux I__9164 (
            .O(N__41316),
            .I(N__41254));
    LocalMux I__9163 (
            .O(N__41307),
            .I(N__41247));
    LocalMux I__9162 (
            .O(N__41302),
            .I(N__41247));
    LocalMux I__9161 (
            .O(N__41293),
            .I(N__41247));
    LocalMux I__9160 (
            .O(N__41284),
            .I(N__41240));
    LocalMux I__9159 (
            .O(N__41275),
            .I(N__41240));
    LocalMux I__9158 (
            .O(N__41266),
            .I(N__41240));
    LocalMux I__9157 (
            .O(N__41257),
            .I(N__41237));
    Span4Mux_h I__9156 (
            .O(N__41254),
            .I(N__41234));
    Span4Mux_v I__9155 (
            .O(N__41247),
            .I(N__41229));
    Span4Mux_v I__9154 (
            .O(N__41240),
            .I(N__41229));
    Span4Mux_h I__9153 (
            .O(N__41237),
            .I(N__41224));
    Span4Mux_h I__9152 (
            .O(N__41234),
            .I(N__41224));
    Odrv4 I__9151 (
            .O(N__41229),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__9150 (
            .O(N__41224),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__9149 (
            .O(N__41219),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CascadeMux I__9148 (
            .O(N__41216),
            .I(N__41213));
    InMux I__9147 (
            .O(N__41213),
            .I(N__41209));
    InMux I__9146 (
            .O(N__41212),
            .I(N__41206));
    LocalMux I__9145 (
            .O(N__41209),
            .I(N__41203));
    LocalMux I__9144 (
            .O(N__41206),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__9143 (
            .O(N__41203),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__9142 (
            .O(N__41198),
            .I(N__41194));
    CEMux I__9141 (
            .O(N__41197),
            .I(N__41190));
    LocalMux I__9140 (
            .O(N__41194),
            .I(N__41187));
    CEMux I__9139 (
            .O(N__41193),
            .I(N__41183));
    LocalMux I__9138 (
            .O(N__41190),
            .I(N__41180));
    Span4Mux_v I__9137 (
            .O(N__41187),
            .I(N__41177));
    CEMux I__9136 (
            .O(N__41186),
            .I(N__41174));
    LocalMux I__9135 (
            .O(N__41183),
            .I(N__41171));
    Span4Mux_v I__9134 (
            .O(N__41180),
            .I(N__41168));
    Span4Mux_h I__9133 (
            .O(N__41177),
            .I(N__41163));
    LocalMux I__9132 (
            .O(N__41174),
            .I(N__41163));
    Span4Mux_h I__9131 (
            .O(N__41171),
            .I(N__41160));
    Span4Mux_h I__9130 (
            .O(N__41168),
            .I(N__41155));
    Span4Mux_h I__9129 (
            .O(N__41163),
            .I(N__41155));
    Odrv4 I__9128 (
            .O(N__41160),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    Odrv4 I__9127 (
            .O(N__41155),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    InMux I__9126 (
            .O(N__41150),
            .I(N__41144));
    InMux I__9125 (
            .O(N__41149),
            .I(N__41141));
    InMux I__9124 (
            .O(N__41148),
            .I(N__41136));
    InMux I__9123 (
            .O(N__41147),
            .I(N__41136));
    LocalMux I__9122 (
            .O(N__41144),
            .I(N__41133));
    LocalMux I__9121 (
            .O(N__41141),
            .I(N__41128));
    LocalMux I__9120 (
            .O(N__41136),
            .I(N__41128));
    Span4Mux_v I__9119 (
            .O(N__41133),
            .I(N__41125));
    Span4Mux_h I__9118 (
            .O(N__41128),
            .I(N__41122));
    Span4Mux_h I__9117 (
            .O(N__41125),
            .I(N__41119));
    Odrv4 I__9116 (
            .O(N__41122),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv4 I__9115 (
            .O(N__41119),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__9114 (
            .O(N__41114),
            .I(N__41106));
    InMux I__9113 (
            .O(N__41113),
            .I(N__41106));
    InMux I__9112 (
            .O(N__41112),
            .I(N__41103));
    InMux I__9111 (
            .O(N__41111),
            .I(N__41100));
    LocalMux I__9110 (
            .O(N__41106),
            .I(N__41097));
    LocalMux I__9109 (
            .O(N__41103),
            .I(N__41094));
    LocalMux I__9108 (
            .O(N__41100),
            .I(N__41091));
    Span4Mux_v I__9107 (
            .O(N__41097),
            .I(N__41088));
    Span4Mux_v I__9106 (
            .O(N__41094),
            .I(N__41085));
    Span4Mux_v I__9105 (
            .O(N__41091),
            .I(N__41082));
    Span4Mux_v I__9104 (
            .O(N__41088),
            .I(N__41079));
    Span4Mux_h I__9103 (
            .O(N__41085),
            .I(N__41076));
    Odrv4 I__9102 (
            .O(N__41082),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv4 I__9101 (
            .O(N__41079),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv4 I__9100 (
            .O(N__41076),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__9099 (
            .O(N__41069),
            .I(N__41066));
    LocalMux I__9098 (
            .O(N__41066),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ));
    InMux I__9097 (
            .O(N__41063),
            .I(N__41059));
    InMux I__9096 (
            .O(N__41062),
            .I(N__41056));
    LocalMux I__9095 (
            .O(N__41059),
            .I(N__41053));
    LocalMux I__9094 (
            .O(N__41056),
            .I(N__41050));
    Span4Mux_h I__9093 (
            .O(N__41053),
            .I(N__41047));
    Span4Mux_v I__9092 (
            .O(N__41050),
            .I(N__41042));
    Span4Mux_h I__9091 (
            .O(N__41047),
            .I(N__41039));
    InMux I__9090 (
            .O(N__41046),
            .I(N__41034));
    InMux I__9089 (
            .O(N__41045),
            .I(N__41034));
    Span4Mux_h I__9088 (
            .O(N__41042),
            .I(N__41031));
    Odrv4 I__9087 (
            .O(N__41039),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    LocalMux I__9086 (
            .O(N__41034),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__9085 (
            .O(N__41031),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__9084 (
            .O(N__41024),
            .I(N__41021));
    LocalMux I__9083 (
            .O(N__41021),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ));
    InMux I__9082 (
            .O(N__41018),
            .I(N__41011));
    InMux I__9081 (
            .O(N__41017),
            .I(N__41011));
    InMux I__9080 (
            .O(N__41016),
            .I(N__41008));
    LocalMux I__9079 (
            .O(N__41011),
            .I(N__41005));
    LocalMux I__9078 (
            .O(N__41008),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv12 I__9077 (
            .O(N__41005),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__9076 (
            .O(N__41000),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    CascadeMux I__9075 (
            .O(N__40997),
            .I(N__40994));
    InMux I__9074 (
            .O(N__40994),
            .I(N__40989));
    InMux I__9073 (
            .O(N__40993),
            .I(N__40986));
    InMux I__9072 (
            .O(N__40992),
            .I(N__40983));
    LocalMux I__9071 (
            .O(N__40989),
            .I(N__40978));
    LocalMux I__9070 (
            .O(N__40986),
            .I(N__40978));
    LocalMux I__9069 (
            .O(N__40983),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv12 I__9068 (
            .O(N__40978),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__9067 (
            .O(N__40973),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__9066 (
            .O(N__40970),
            .I(N__40966));
    CascadeMux I__9065 (
            .O(N__40969),
            .I(N__40963));
    InMux I__9064 (
            .O(N__40966),
            .I(N__40957));
    InMux I__9063 (
            .O(N__40963),
            .I(N__40957));
    InMux I__9062 (
            .O(N__40962),
            .I(N__40954));
    LocalMux I__9061 (
            .O(N__40957),
            .I(N__40951));
    LocalMux I__9060 (
            .O(N__40954),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__9059 (
            .O(N__40951),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__9058 (
            .O(N__40946),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__9057 (
            .O(N__40943),
            .I(N__40936));
    InMux I__9056 (
            .O(N__40942),
            .I(N__40936));
    InMux I__9055 (
            .O(N__40941),
            .I(N__40933));
    LocalMux I__9054 (
            .O(N__40936),
            .I(N__40930));
    LocalMux I__9053 (
            .O(N__40933),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv12 I__9052 (
            .O(N__40930),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__9051 (
            .O(N__40925),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__9050 (
            .O(N__40922),
            .I(N__40915));
    InMux I__9049 (
            .O(N__40921),
            .I(N__40915));
    InMux I__9048 (
            .O(N__40920),
            .I(N__40912));
    LocalMux I__9047 (
            .O(N__40915),
            .I(N__40909));
    LocalMux I__9046 (
            .O(N__40912),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__9045 (
            .O(N__40909),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__9044 (
            .O(N__40904),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__9043 (
            .O(N__40901),
            .I(N__40897));
    CascadeMux I__9042 (
            .O(N__40900),
            .I(N__40894));
    InMux I__9041 (
            .O(N__40897),
            .I(N__40888));
    InMux I__9040 (
            .O(N__40894),
            .I(N__40888));
    InMux I__9039 (
            .O(N__40893),
            .I(N__40885));
    LocalMux I__9038 (
            .O(N__40888),
            .I(N__40882));
    LocalMux I__9037 (
            .O(N__40885),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__9036 (
            .O(N__40882),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__9035 (
            .O(N__40877),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__9034 (
            .O(N__40874),
            .I(N__40870));
    CascadeMux I__9033 (
            .O(N__40873),
            .I(N__40867));
    InMux I__9032 (
            .O(N__40870),
            .I(N__40864));
    InMux I__9031 (
            .O(N__40867),
            .I(N__40860));
    LocalMux I__9030 (
            .O(N__40864),
            .I(N__40857));
    InMux I__9029 (
            .O(N__40863),
            .I(N__40854));
    LocalMux I__9028 (
            .O(N__40860),
            .I(N__40851));
    Span4Mux_v I__9027 (
            .O(N__40857),
            .I(N__40848));
    LocalMux I__9026 (
            .O(N__40854),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv12 I__9025 (
            .O(N__40851),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv4 I__9024 (
            .O(N__40848),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__9023 (
            .O(N__40841),
            .I(bfn_17_21_0_));
    CascadeMux I__9022 (
            .O(N__40838),
            .I(N__40834));
    InMux I__9021 (
            .O(N__40837),
            .I(N__40831));
    InMux I__9020 (
            .O(N__40834),
            .I(N__40827));
    LocalMux I__9019 (
            .O(N__40831),
            .I(N__40824));
    InMux I__9018 (
            .O(N__40830),
            .I(N__40821));
    LocalMux I__9017 (
            .O(N__40827),
            .I(N__40818));
    Span4Mux_v I__9016 (
            .O(N__40824),
            .I(N__40815));
    LocalMux I__9015 (
            .O(N__40821),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv12 I__9014 (
            .O(N__40818),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__9013 (
            .O(N__40815),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__9012 (
            .O(N__40808),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__9011 (
            .O(N__40805),
            .I(N__40798));
    InMux I__9010 (
            .O(N__40804),
            .I(N__40798));
    InMux I__9009 (
            .O(N__40803),
            .I(N__40795));
    LocalMux I__9008 (
            .O(N__40798),
            .I(N__40792));
    LocalMux I__9007 (
            .O(N__40795),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__9006 (
            .O(N__40792),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__9005 (
            .O(N__40787),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__9004 (
            .O(N__40784),
            .I(N__40777));
    InMux I__9003 (
            .O(N__40783),
            .I(N__40777));
    InMux I__9002 (
            .O(N__40782),
            .I(N__40774));
    LocalMux I__9001 (
            .O(N__40777),
            .I(N__40771));
    LocalMux I__9000 (
            .O(N__40774),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__8999 (
            .O(N__40771),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__8998 (
            .O(N__40766),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__8997 (
            .O(N__40763),
            .I(N__40756));
    InMux I__8996 (
            .O(N__40762),
            .I(N__40756));
    InMux I__8995 (
            .O(N__40761),
            .I(N__40753));
    LocalMux I__8994 (
            .O(N__40756),
            .I(N__40750));
    LocalMux I__8993 (
            .O(N__40753),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__8992 (
            .O(N__40750),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__8991 (
            .O(N__40745),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__8990 (
            .O(N__40742),
            .I(N__40738));
    InMux I__8989 (
            .O(N__40741),
            .I(N__40734));
    InMux I__8988 (
            .O(N__40738),
            .I(N__40731));
    InMux I__8987 (
            .O(N__40737),
            .I(N__40728));
    LocalMux I__8986 (
            .O(N__40734),
            .I(N__40723));
    LocalMux I__8985 (
            .O(N__40731),
            .I(N__40723));
    LocalMux I__8984 (
            .O(N__40728),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__8983 (
            .O(N__40723),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__8982 (
            .O(N__40718),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__8981 (
            .O(N__40715),
            .I(N__40711));
    InMux I__8980 (
            .O(N__40714),
            .I(N__40707));
    InMux I__8979 (
            .O(N__40711),
            .I(N__40704));
    InMux I__8978 (
            .O(N__40710),
            .I(N__40701));
    LocalMux I__8977 (
            .O(N__40707),
            .I(N__40696));
    LocalMux I__8976 (
            .O(N__40704),
            .I(N__40696));
    LocalMux I__8975 (
            .O(N__40701),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__8974 (
            .O(N__40696),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__8973 (
            .O(N__40691),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__8972 (
            .O(N__40688),
            .I(N__40684));
    CascadeMux I__8971 (
            .O(N__40687),
            .I(N__40681));
    InMux I__8970 (
            .O(N__40684),
            .I(N__40675));
    InMux I__8969 (
            .O(N__40681),
            .I(N__40675));
    InMux I__8968 (
            .O(N__40680),
            .I(N__40672));
    LocalMux I__8967 (
            .O(N__40675),
            .I(N__40669));
    LocalMux I__8966 (
            .O(N__40672),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__8965 (
            .O(N__40669),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__8964 (
            .O(N__40664),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    CascadeMux I__8963 (
            .O(N__40661),
            .I(N__40657));
    CascadeMux I__8962 (
            .O(N__40660),
            .I(N__40654));
    InMux I__8961 (
            .O(N__40657),
            .I(N__40648));
    InMux I__8960 (
            .O(N__40654),
            .I(N__40648));
    InMux I__8959 (
            .O(N__40653),
            .I(N__40645));
    LocalMux I__8958 (
            .O(N__40648),
            .I(N__40642));
    LocalMux I__8957 (
            .O(N__40645),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__8956 (
            .O(N__40642),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__8955 (
            .O(N__40637),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__8954 (
            .O(N__40634),
            .I(N__40630));
    InMux I__8953 (
            .O(N__40633),
            .I(N__40627));
    InMux I__8952 (
            .O(N__40630),
            .I(N__40623));
    LocalMux I__8951 (
            .O(N__40627),
            .I(N__40620));
    InMux I__8950 (
            .O(N__40626),
            .I(N__40617));
    LocalMux I__8949 (
            .O(N__40623),
            .I(N__40614));
    Span4Mux_v I__8948 (
            .O(N__40620),
            .I(N__40611));
    LocalMux I__8947 (
            .O(N__40617),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv12 I__8946 (
            .O(N__40614),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv4 I__8945 (
            .O(N__40611),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__8944 (
            .O(N__40604),
            .I(bfn_17_20_0_));
    CascadeMux I__8943 (
            .O(N__40601),
            .I(N__40597));
    InMux I__8942 (
            .O(N__40600),
            .I(N__40594));
    InMux I__8941 (
            .O(N__40597),
            .I(N__40591));
    LocalMux I__8940 (
            .O(N__40594),
            .I(N__40588));
    LocalMux I__8939 (
            .O(N__40591),
            .I(N__40582));
    Span4Mux_v I__8938 (
            .O(N__40588),
            .I(N__40582));
    InMux I__8937 (
            .O(N__40587),
            .I(N__40579));
    Span4Mux_h I__8936 (
            .O(N__40582),
            .I(N__40576));
    LocalMux I__8935 (
            .O(N__40579),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__8934 (
            .O(N__40576),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__8933 (
            .O(N__40571),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__8932 (
            .O(N__40568),
            .I(N__40561));
    InMux I__8931 (
            .O(N__40567),
            .I(N__40561));
    InMux I__8930 (
            .O(N__40566),
            .I(N__40558));
    LocalMux I__8929 (
            .O(N__40561),
            .I(N__40555));
    LocalMux I__8928 (
            .O(N__40558),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__8927 (
            .O(N__40555),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__8926 (
            .O(N__40550),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    CascadeMux I__8925 (
            .O(N__40547),
            .I(N__40543));
    InMux I__8924 (
            .O(N__40546),
            .I(N__40540));
    InMux I__8923 (
            .O(N__40543),
            .I(N__40537));
    LocalMux I__8922 (
            .O(N__40540),
            .I(N__40531));
    LocalMux I__8921 (
            .O(N__40537),
            .I(N__40531));
    InMux I__8920 (
            .O(N__40536),
            .I(N__40528));
    Span4Mux_h I__8919 (
            .O(N__40531),
            .I(N__40525));
    LocalMux I__8918 (
            .O(N__40528),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__8917 (
            .O(N__40525),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__8916 (
            .O(N__40520),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__8915 (
            .O(N__40517),
            .I(N__40513));
    CascadeMux I__8914 (
            .O(N__40516),
            .I(N__40510));
    InMux I__8913 (
            .O(N__40513),
            .I(N__40504));
    InMux I__8912 (
            .O(N__40510),
            .I(N__40504));
    InMux I__8911 (
            .O(N__40509),
            .I(N__40501));
    LocalMux I__8910 (
            .O(N__40504),
            .I(N__40498));
    LocalMux I__8909 (
            .O(N__40501),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__8908 (
            .O(N__40498),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__8907 (
            .O(N__40493),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__8906 (
            .O(N__40490),
            .I(N__40486));
    CascadeMux I__8905 (
            .O(N__40489),
            .I(N__40483));
    InMux I__8904 (
            .O(N__40486),
            .I(N__40477));
    InMux I__8903 (
            .O(N__40483),
            .I(N__40477));
    InMux I__8902 (
            .O(N__40482),
            .I(N__40474));
    LocalMux I__8901 (
            .O(N__40477),
            .I(N__40471));
    LocalMux I__8900 (
            .O(N__40474),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__8899 (
            .O(N__40471),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__8898 (
            .O(N__40466),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__8897 (
            .O(N__40463),
            .I(N__40456));
    InMux I__8896 (
            .O(N__40462),
            .I(N__40456));
    InMux I__8895 (
            .O(N__40461),
            .I(N__40453));
    LocalMux I__8894 (
            .O(N__40456),
            .I(N__40450));
    LocalMux I__8893 (
            .O(N__40453),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__8892 (
            .O(N__40450),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__8891 (
            .O(N__40445),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__8890 (
            .O(N__40442),
            .I(N__40435));
    InMux I__8889 (
            .O(N__40441),
            .I(N__40435));
    InMux I__8888 (
            .O(N__40440),
            .I(N__40432));
    LocalMux I__8887 (
            .O(N__40435),
            .I(N__40429));
    LocalMux I__8886 (
            .O(N__40432),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__8885 (
            .O(N__40429),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__8884 (
            .O(N__40424),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__8883 (
            .O(N__40421),
            .I(N__40417));
    CascadeMux I__8882 (
            .O(N__40420),
            .I(N__40414));
    InMux I__8881 (
            .O(N__40417),
            .I(N__40410));
    InMux I__8880 (
            .O(N__40414),
            .I(N__40407));
    InMux I__8879 (
            .O(N__40413),
            .I(N__40404));
    LocalMux I__8878 (
            .O(N__40410),
            .I(N__40399));
    LocalMux I__8877 (
            .O(N__40407),
            .I(N__40399));
    LocalMux I__8876 (
            .O(N__40404),
            .I(N__40394));
    Span4Mux_v I__8875 (
            .O(N__40399),
            .I(N__40394));
    Odrv4 I__8874 (
            .O(N__40394),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__8873 (
            .O(N__40391),
            .I(bfn_17_19_0_));
    CascadeMux I__8872 (
            .O(N__40388),
            .I(N__40384));
    CascadeMux I__8871 (
            .O(N__40387),
            .I(N__40381));
    InMux I__8870 (
            .O(N__40384),
            .I(N__40378));
    InMux I__8869 (
            .O(N__40381),
            .I(N__40375));
    LocalMux I__8868 (
            .O(N__40378),
            .I(N__40371));
    LocalMux I__8867 (
            .O(N__40375),
            .I(N__40368));
    InMux I__8866 (
            .O(N__40374),
            .I(N__40365));
    Span4Mux_h I__8865 (
            .O(N__40371),
            .I(N__40360));
    Span4Mux_v I__8864 (
            .O(N__40368),
            .I(N__40360));
    LocalMux I__8863 (
            .O(N__40365),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__8862 (
            .O(N__40360),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__8861 (
            .O(N__40355),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    CascadeMux I__8860 (
            .O(N__40352),
            .I(N__40349));
    InMux I__8859 (
            .O(N__40349),
            .I(N__40344));
    InMux I__8858 (
            .O(N__40348),
            .I(N__40341));
    InMux I__8857 (
            .O(N__40347),
            .I(N__40338));
    LocalMux I__8856 (
            .O(N__40344),
            .I(N__40335));
    LocalMux I__8855 (
            .O(N__40341),
            .I(N__40332));
    LocalMux I__8854 (
            .O(N__40338),
            .I(N__40329));
    Span4Mux_v I__8853 (
            .O(N__40335),
            .I(N__40323));
    Span4Mux_h I__8852 (
            .O(N__40332),
            .I(N__40323));
    Span4Mux_h I__8851 (
            .O(N__40329),
            .I(N__40320));
    InMux I__8850 (
            .O(N__40328),
            .I(N__40317));
    Odrv4 I__8849 (
            .O(N__40323),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__8848 (
            .O(N__40320),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__8847 (
            .O(N__40317),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__8846 (
            .O(N__40310),
            .I(N__40307));
    LocalMux I__8845 (
            .O(N__40307),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__8844 (
            .O(N__40304),
            .I(N__40297));
    InMux I__8843 (
            .O(N__40303),
            .I(N__40297));
    InMux I__8842 (
            .O(N__40302),
            .I(N__40294));
    LocalMux I__8841 (
            .O(N__40297),
            .I(N__40289));
    LocalMux I__8840 (
            .O(N__40294),
            .I(N__40289));
    Span4Mux_h I__8839 (
            .O(N__40289),
            .I(N__40285));
    InMux I__8838 (
            .O(N__40288),
            .I(N__40282));
    Odrv4 I__8837 (
            .O(N__40285),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__8836 (
            .O(N__40282),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    CascadeMux I__8835 (
            .O(N__40277),
            .I(N__40274));
    InMux I__8834 (
            .O(N__40274),
            .I(N__40271));
    LocalMux I__8833 (
            .O(N__40271),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__8832 (
            .O(N__40268),
            .I(N__40265));
    LocalMux I__8831 (
            .O(N__40265),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__8830 (
            .O(N__40262),
            .I(N__40255));
    InMux I__8829 (
            .O(N__40261),
            .I(N__40255));
    InMux I__8828 (
            .O(N__40260),
            .I(N__40252));
    LocalMux I__8827 (
            .O(N__40255),
            .I(N__40249));
    LocalMux I__8826 (
            .O(N__40252),
            .I(N__40245));
    Span4Mux_h I__8825 (
            .O(N__40249),
            .I(N__40242));
    InMux I__8824 (
            .O(N__40248),
            .I(N__40239));
    Odrv12 I__8823 (
            .O(N__40245),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    Odrv4 I__8822 (
            .O(N__40242),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__8821 (
            .O(N__40239),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    CascadeMux I__8820 (
            .O(N__40232),
            .I(N__40229));
    InMux I__8819 (
            .O(N__40229),
            .I(N__40226));
    LocalMux I__8818 (
            .O(N__40226),
            .I(N__40223));
    Span4Mux_v I__8817 (
            .O(N__40223),
            .I(N__40220));
    Span4Mux_h I__8816 (
            .O(N__40220),
            .I(N__40217));
    Odrv4 I__8815 (
            .O(N__40217),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__8814 (
            .O(N__40214),
            .I(N__40211));
    LocalMux I__8813 (
            .O(N__40211),
            .I(N__40208));
    Odrv12 I__8812 (
            .O(N__40208),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__8811 (
            .O(N__40205),
            .I(N__40202));
    LocalMux I__8810 (
            .O(N__40202),
            .I(N__40199));
    Span4Mux_h I__8809 (
            .O(N__40199),
            .I(N__40196));
    Odrv4 I__8808 (
            .O(N__40196),
            .I(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ));
    InMux I__8807 (
            .O(N__40193),
            .I(N__40188));
    InMux I__8806 (
            .O(N__40192),
            .I(N__40185));
    InMux I__8805 (
            .O(N__40191),
            .I(N__40182));
    LocalMux I__8804 (
            .O(N__40188),
            .I(N__40179));
    LocalMux I__8803 (
            .O(N__40185),
            .I(N__40175));
    LocalMux I__8802 (
            .O(N__40182),
            .I(N__40170));
    Span4Mux_h I__8801 (
            .O(N__40179),
            .I(N__40170));
    InMux I__8800 (
            .O(N__40178),
            .I(N__40167));
    Odrv12 I__8799 (
            .O(N__40175),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    Odrv4 I__8798 (
            .O(N__40170),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__8797 (
            .O(N__40167),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__8796 (
            .O(N__40160),
            .I(N__40157));
    LocalMux I__8795 (
            .O(N__40157),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__8794 (
            .O(N__40154),
            .I(N__40150));
    CascadeMux I__8793 (
            .O(N__40153),
            .I(N__40147));
    LocalMux I__8792 (
            .O(N__40150),
            .I(N__40143));
    InMux I__8791 (
            .O(N__40147),
            .I(N__40140));
    InMux I__8790 (
            .O(N__40146),
            .I(N__40137));
    Span12Mux_v I__8789 (
            .O(N__40143),
            .I(N__40132));
    LocalMux I__8788 (
            .O(N__40140),
            .I(N__40132));
    LocalMux I__8787 (
            .O(N__40137),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv12 I__8786 (
            .O(N__40132),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__8785 (
            .O(N__40127),
            .I(bfn_17_18_0_));
    InMux I__8784 (
            .O(N__40124),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    CascadeMux I__8783 (
            .O(N__40121),
            .I(N__40117));
    InMux I__8782 (
            .O(N__40120),
            .I(N__40114));
    InMux I__8781 (
            .O(N__40117),
            .I(N__40110));
    LocalMux I__8780 (
            .O(N__40114),
            .I(N__40107));
    InMux I__8779 (
            .O(N__40113),
            .I(N__40104));
    LocalMux I__8778 (
            .O(N__40110),
            .I(N__40101));
    Span4Mux_v I__8777 (
            .O(N__40107),
            .I(N__40096));
    LocalMux I__8776 (
            .O(N__40104),
            .I(N__40096));
    Span4Mux_h I__8775 (
            .O(N__40101),
            .I(N__40090));
    Span4Mux_h I__8774 (
            .O(N__40096),
            .I(N__40090));
    InMux I__8773 (
            .O(N__40095),
            .I(N__40087));
    Odrv4 I__8772 (
            .O(N__40090),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__8771 (
            .O(N__40087),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    CascadeMux I__8770 (
            .O(N__40082),
            .I(N__40079));
    InMux I__8769 (
            .O(N__40079),
            .I(N__40076));
    LocalMux I__8768 (
            .O(N__40076),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    InMux I__8767 (
            .O(N__40073),
            .I(N__40069));
    InMux I__8766 (
            .O(N__40072),
            .I(N__40066));
    LocalMux I__8765 (
            .O(N__40069),
            .I(N__40062));
    LocalMux I__8764 (
            .O(N__40066),
            .I(N__40059));
    InMux I__8763 (
            .O(N__40065),
            .I(N__40056));
    Span4Mux_h I__8762 (
            .O(N__40062),
            .I(N__40053));
    Span4Mux_h I__8761 (
            .O(N__40059),
            .I(N__40049));
    LocalMux I__8760 (
            .O(N__40056),
            .I(N__40046));
    Span4Mux_v I__8759 (
            .O(N__40053),
            .I(N__40043));
    InMux I__8758 (
            .O(N__40052),
            .I(N__40040));
    Odrv4 I__8757 (
            .O(N__40049),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv12 I__8756 (
            .O(N__40046),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__8755 (
            .O(N__40043),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__8754 (
            .O(N__40040),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    CascadeMux I__8753 (
            .O(N__40031),
            .I(N__40028));
    InMux I__8752 (
            .O(N__40028),
            .I(N__40025));
    LocalMux I__8751 (
            .O(N__40025),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    InMux I__8750 (
            .O(N__40022),
            .I(N__40019));
    LocalMux I__8749 (
            .O(N__40019),
            .I(N__40014));
    InMux I__8748 (
            .O(N__40018),
            .I(N__40011));
    InMux I__8747 (
            .O(N__40017),
            .I(N__40008));
    Span4Mux_v I__8746 (
            .O(N__40014),
            .I(N__40003));
    LocalMux I__8745 (
            .O(N__40011),
            .I(N__40003));
    LocalMux I__8744 (
            .O(N__40008),
            .I(N__40000));
    Span4Mux_h I__8743 (
            .O(N__40003),
            .I(N__39994));
    Span4Mux_h I__8742 (
            .O(N__40000),
            .I(N__39994));
    InMux I__8741 (
            .O(N__39999),
            .I(N__39991));
    Odrv4 I__8740 (
            .O(N__39994),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__8739 (
            .O(N__39991),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    CascadeMux I__8738 (
            .O(N__39986),
            .I(N__39983));
    InMux I__8737 (
            .O(N__39983),
            .I(N__39980));
    LocalMux I__8736 (
            .O(N__39980),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__8735 (
            .O(N__39977),
            .I(N__39974));
    LocalMux I__8734 (
            .O(N__39974),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    InMux I__8733 (
            .O(N__39971),
            .I(N__39966));
    InMux I__8732 (
            .O(N__39970),
            .I(N__39963));
    InMux I__8731 (
            .O(N__39969),
            .I(N__39960));
    LocalMux I__8730 (
            .O(N__39966),
            .I(N__39957));
    LocalMux I__8729 (
            .O(N__39963),
            .I(N__39952));
    LocalMux I__8728 (
            .O(N__39960),
            .I(N__39952));
    Span4Mux_h I__8727 (
            .O(N__39957),
            .I(N__39946));
    Span4Mux_h I__8726 (
            .O(N__39952),
            .I(N__39946));
    InMux I__8725 (
            .O(N__39951),
            .I(N__39943));
    Odrv4 I__8724 (
            .O(N__39946),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__8723 (
            .O(N__39943),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__8722 (
            .O(N__39938),
            .I(N__39935));
    LocalMux I__8721 (
            .O(N__39935),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__8720 (
            .O(N__39932),
            .I(N__39929));
    LocalMux I__8719 (
            .O(N__39929),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__8718 (
            .O(N__39926),
            .I(N__39922));
    CascadeMux I__8717 (
            .O(N__39925),
            .I(N__39919));
    InMux I__8716 (
            .O(N__39922),
            .I(N__39915));
    InMux I__8715 (
            .O(N__39919),
            .I(N__39912));
    InMux I__8714 (
            .O(N__39918),
            .I(N__39909));
    LocalMux I__8713 (
            .O(N__39915),
            .I(N__39904));
    LocalMux I__8712 (
            .O(N__39912),
            .I(N__39904));
    LocalMux I__8711 (
            .O(N__39909),
            .I(N__39901));
    Span4Mux_h I__8710 (
            .O(N__39904),
            .I(N__39895));
    Span4Mux_h I__8709 (
            .O(N__39901),
            .I(N__39895));
    InMux I__8708 (
            .O(N__39900),
            .I(N__39892));
    Odrv4 I__8707 (
            .O(N__39895),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__8706 (
            .O(N__39892),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    CascadeMux I__8705 (
            .O(N__39887),
            .I(N__39884));
    InMux I__8704 (
            .O(N__39884),
            .I(N__39881));
    LocalMux I__8703 (
            .O(N__39881),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__8702 (
            .O(N__39878),
            .I(N__39873));
    InMux I__8701 (
            .O(N__39877),
            .I(N__39870));
    InMux I__8700 (
            .O(N__39876),
            .I(N__39867));
    LocalMux I__8699 (
            .O(N__39873),
            .I(N__39864));
    LocalMux I__8698 (
            .O(N__39870),
            .I(N__39861));
    LocalMux I__8697 (
            .O(N__39867),
            .I(N__39857));
    Span4Mux_h I__8696 (
            .O(N__39864),
            .I(N__39852));
    Span4Mux_h I__8695 (
            .O(N__39861),
            .I(N__39852));
    InMux I__8694 (
            .O(N__39860),
            .I(N__39849));
    Odrv12 I__8693 (
            .O(N__39857),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    Odrv4 I__8692 (
            .O(N__39852),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__8691 (
            .O(N__39849),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    CascadeMux I__8690 (
            .O(N__39842),
            .I(N__39839));
    InMux I__8689 (
            .O(N__39839),
            .I(N__39836));
    LocalMux I__8688 (
            .O(N__39836),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    CascadeMux I__8687 (
            .O(N__39833),
            .I(N__39830));
    InMux I__8686 (
            .O(N__39830),
            .I(N__39827));
    LocalMux I__8685 (
            .O(N__39827),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    CascadeMux I__8684 (
            .O(N__39824),
            .I(N__39819));
    CascadeMux I__8683 (
            .O(N__39823),
            .I(N__39816));
    InMux I__8682 (
            .O(N__39822),
            .I(N__39813));
    InMux I__8681 (
            .O(N__39819),
            .I(N__39808));
    InMux I__8680 (
            .O(N__39816),
            .I(N__39808));
    LocalMux I__8679 (
            .O(N__39813),
            .I(N__39805));
    LocalMux I__8678 (
            .O(N__39808),
            .I(N__39801));
    Span4Mux_h I__8677 (
            .O(N__39805),
            .I(N__39798));
    InMux I__8676 (
            .O(N__39804),
            .I(N__39795));
    Odrv12 I__8675 (
            .O(N__39801),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__8674 (
            .O(N__39798),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__8673 (
            .O(N__39795),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    CascadeMux I__8672 (
            .O(N__39788),
            .I(N__39785));
    InMux I__8671 (
            .O(N__39785),
            .I(N__39782));
    LocalMux I__8670 (
            .O(N__39782),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    CascadeMux I__8669 (
            .O(N__39779),
            .I(N__39776));
    InMux I__8668 (
            .O(N__39776),
            .I(N__39773));
    LocalMux I__8667 (
            .O(N__39773),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    CascadeMux I__8666 (
            .O(N__39770),
            .I(N__39767));
    InMux I__8665 (
            .O(N__39767),
            .I(N__39764));
    LocalMux I__8664 (
            .O(N__39764),
            .I(N__39761));
    Odrv12 I__8663 (
            .O(N__39761),
            .I(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ));
    CascadeMux I__8662 (
            .O(N__39758),
            .I(N__39754));
    CascadeMux I__8661 (
            .O(N__39757),
            .I(N__39751));
    InMux I__8660 (
            .O(N__39754),
            .I(N__39747));
    InMux I__8659 (
            .O(N__39751),
            .I(N__39744));
    InMux I__8658 (
            .O(N__39750),
            .I(N__39741));
    LocalMux I__8657 (
            .O(N__39747),
            .I(N__39736));
    LocalMux I__8656 (
            .O(N__39744),
            .I(N__39736));
    LocalMux I__8655 (
            .O(N__39741),
            .I(N__39733));
    Span4Mux_h I__8654 (
            .O(N__39736),
            .I(N__39728));
    Span4Mux_h I__8653 (
            .O(N__39733),
            .I(N__39728));
    Span4Mux_v I__8652 (
            .O(N__39728),
            .I(N__39724));
    InMux I__8651 (
            .O(N__39727),
            .I(N__39721));
    Odrv4 I__8650 (
            .O(N__39724),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__8649 (
            .O(N__39721),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__8648 (
            .O(N__39716),
            .I(N__39713));
    LocalMux I__8647 (
            .O(N__39713),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__8646 (
            .O(N__39710),
            .I(N__39706));
    CascadeMux I__8645 (
            .O(N__39709),
            .I(N__39703));
    InMux I__8644 (
            .O(N__39706),
            .I(N__39697));
    InMux I__8643 (
            .O(N__39703),
            .I(N__39697));
    InMux I__8642 (
            .O(N__39702),
            .I(N__39694));
    LocalMux I__8641 (
            .O(N__39697),
            .I(N__39691));
    LocalMux I__8640 (
            .O(N__39694),
            .I(N__39688));
    Span4Mux_h I__8639 (
            .O(N__39691),
            .I(N__39682));
    Span4Mux_h I__8638 (
            .O(N__39688),
            .I(N__39682));
    InMux I__8637 (
            .O(N__39687),
            .I(N__39679));
    Odrv4 I__8636 (
            .O(N__39682),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__8635 (
            .O(N__39679),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    CascadeMux I__8634 (
            .O(N__39674),
            .I(N__39671));
    InMux I__8633 (
            .O(N__39671),
            .I(N__39668));
    LocalMux I__8632 (
            .O(N__39668),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    CascadeMux I__8631 (
            .O(N__39665),
            .I(N__39661));
    InMux I__8630 (
            .O(N__39664),
            .I(N__39657));
    InMux I__8629 (
            .O(N__39661),
            .I(N__39654));
    InMux I__8628 (
            .O(N__39660),
            .I(N__39651));
    LocalMux I__8627 (
            .O(N__39657),
            .I(N__39648));
    LocalMux I__8626 (
            .O(N__39654),
            .I(N__39643));
    LocalMux I__8625 (
            .O(N__39651),
            .I(N__39643));
    Span4Mux_h I__8624 (
            .O(N__39648),
            .I(N__39637));
    Span4Mux_h I__8623 (
            .O(N__39643),
            .I(N__39637));
    InMux I__8622 (
            .O(N__39642),
            .I(N__39634));
    Odrv4 I__8621 (
            .O(N__39637),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__8620 (
            .O(N__39634),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    CascadeMux I__8619 (
            .O(N__39629),
            .I(N__39626));
    InMux I__8618 (
            .O(N__39626),
            .I(N__39623));
    LocalMux I__8617 (
            .O(N__39623),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    CascadeMux I__8616 (
            .O(N__39620),
            .I(N__39616));
    CascadeMux I__8615 (
            .O(N__39619),
            .I(N__39612));
    InMux I__8614 (
            .O(N__39616),
            .I(N__39609));
    InMux I__8613 (
            .O(N__39615),
            .I(N__39606));
    InMux I__8612 (
            .O(N__39612),
            .I(N__39603));
    LocalMux I__8611 (
            .O(N__39609),
            .I(N__39600));
    LocalMux I__8610 (
            .O(N__39606),
            .I(N__39597));
    LocalMux I__8609 (
            .O(N__39603),
            .I(N__39593));
    Span4Mux_h I__8608 (
            .O(N__39600),
            .I(N__39588));
    Span4Mux_h I__8607 (
            .O(N__39597),
            .I(N__39588));
    InMux I__8606 (
            .O(N__39596),
            .I(N__39585));
    Odrv12 I__8605 (
            .O(N__39593),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__8604 (
            .O(N__39588),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__8603 (
            .O(N__39585),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__8602 (
            .O(N__39578),
            .I(N__39575));
    LocalMux I__8601 (
            .O(N__39575),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    InMux I__8600 (
            .O(N__39572),
            .I(N__39568));
    InMux I__8599 (
            .O(N__39571),
            .I(N__39564));
    LocalMux I__8598 (
            .O(N__39568),
            .I(N__39561));
    InMux I__8597 (
            .O(N__39567),
            .I(N__39558));
    LocalMux I__8596 (
            .O(N__39564),
            .I(N__39553));
    Span4Mux_h I__8595 (
            .O(N__39561),
            .I(N__39553));
    LocalMux I__8594 (
            .O(N__39558),
            .I(N__39549));
    Span4Mux_h I__8593 (
            .O(N__39553),
            .I(N__39546));
    InMux I__8592 (
            .O(N__39552),
            .I(N__39543));
    Odrv12 I__8591 (
            .O(N__39549),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__8590 (
            .O(N__39546),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__8589 (
            .O(N__39543),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    InMux I__8588 (
            .O(N__39536),
            .I(N__39533));
    LocalMux I__8587 (
            .O(N__39533),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    InMux I__8586 (
            .O(N__39530),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    CascadeMux I__8585 (
            .O(N__39527),
            .I(N__39522));
    InMux I__8584 (
            .O(N__39526),
            .I(N__39517));
    InMux I__8583 (
            .O(N__39525),
            .I(N__39517));
    InMux I__8582 (
            .O(N__39522),
            .I(N__39513));
    LocalMux I__8581 (
            .O(N__39517),
            .I(N__39510));
    InMux I__8580 (
            .O(N__39516),
            .I(N__39507));
    LocalMux I__8579 (
            .O(N__39513),
            .I(N__39504));
    Span4Mux_h I__8578 (
            .O(N__39510),
            .I(N__39501));
    LocalMux I__8577 (
            .O(N__39507),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv12 I__8576 (
            .O(N__39504),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__8575 (
            .O(N__39501),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__8574 (
            .O(N__39494),
            .I(N__39490));
    InMux I__8573 (
            .O(N__39493),
            .I(N__39486));
    LocalMux I__8572 (
            .O(N__39490),
            .I(N__39483));
    InMux I__8571 (
            .O(N__39489),
            .I(N__39480));
    LocalMux I__8570 (
            .O(N__39486),
            .I(N__39475));
    Span4Mux_h I__8569 (
            .O(N__39483),
            .I(N__39475));
    LocalMux I__8568 (
            .O(N__39480),
            .I(N__39471));
    Span4Mux_v I__8567 (
            .O(N__39475),
            .I(N__39468));
    InMux I__8566 (
            .O(N__39474),
            .I(N__39465));
    Odrv12 I__8565 (
            .O(N__39471),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    Odrv4 I__8564 (
            .O(N__39468),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__8563 (
            .O(N__39465),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__8562 (
            .O(N__39458),
            .I(N__39455));
    LocalMux I__8561 (
            .O(N__39455),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__8560 (
            .O(N__39452),
            .I(N__39449));
    LocalMux I__8559 (
            .O(N__39449),
            .I(N__39444));
    InMux I__8558 (
            .O(N__39448),
            .I(N__39441));
    InMux I__8557 (
            .O(N__39447),
            .I(N__39438));
    Span4Mux_h I__8556 (
            .O(N__39444),
            .I(N__39435));
    LocalMux I__8555 (
            .O(N__39441),
            .I(N__39429));
    LocalMux I__8554 (
            .O(N__39438),
            .I(N__39429));
    Span4Mux_v I__8553 (
            .O(N__39435),
            .I(N__39426));
    InMux I__8552 (
            .O(N__39434),
            .I(N__39423));
    Odrv12 I__8551 (
            .O(N__39429),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__8550 (
            .O(N__39426),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__8549 (
            .O(N__39423),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    CascadeMux I__8548 (
            .O(N__39416),
            .I(N__39413));
    InMux I__8547 (
            .O(N__39413),
            .I(N__39410));
    LocalMux I__8546 (
            .O(N__39410),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__8545 (
            .O(N__39407),
            .I(N__39400));
    InMux I__8544 (
            .O(N__39406),
            .I(N__39400));
    InMux I__8543 (
            .O(N__39405),
            .I(N__39397));
    LocalMux I__8542 (
            .O(N__39400),
            .I(N__39392));
    LocalMux I__8541 (
            .O(N__39397),
            .I(N__39392));
    Span4Mux_h I__8540 (
            .O(N__39392),
            .I(N__39388));
    InMux I__8539 (
            .O(N__39391),
            .I(N__39385));
    Odrv4 I__8538 (
            .O(N__39388),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__8537 (
            .O(N__39385),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__8536 (
            .O(N__39380),
            .I(N__39377));
    LocalMux I__8535 (
            .O(N__39377),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__8534 (
            .O(N__39374),
            .I(N__39370));
    CascadeMux I__8533 (
            .O(N__39373),
            .I(N__39366));
    InMux I__8532 (
            .O(N__39370),
            .I(N__39363));
    InMux I__8531 (
            .O(N__39369),
            .I(N__39360));
    InMux I__8530 (
            .O(N__39366),
            .I(N__39357));
    LocalMux I__8529 (
            .O(N__39363),
            .I(N__39354));
    LocalMux I__8528 (
            .O(N__39360),
            .I(N__39351));
    LocalMux I__8527 (
            .O(N__39357),
            .I(N__39343));
    Span4Mux_h I__8526 (
            .O(N__39354),
            .I(N__39343));
    Span4Mux_h I__8525 (
            .O(N__39351),
            .I(N__39343));
    InMux I__8524 (
            .O(N__39350),
            .I(N__39340));
    Odrv4 I__8523 (
            .O(N__39343),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__8522 (
            .O(N__39340),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    CascadeMux I__8521 (
            .O(N__39335),
            .I(N__39332));
    InMux I__8520 (
            .O(N__39332),
            .I(N__39329));
    LocalMux I__8519 (
            .O(N__39329),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__8518 (
            .O(N__39326),
            .I(N__39322));
    InMux I__8517 (
            .O(N__39325),
            .I(N__39316));
    InMux I__8516 (
            .O(N__39322),
            .I(N__39316));
    InMux I__8515 (
            .O(N__39321),
            .I(N__39313));
    LocalMux I__8514 (
            .O(N__39316),
            .I(N__39310));
    LocalMux I__8513 (
            .O(N__39313),
            .I(N__39307));
    Span4Mux_h I__8512 (
            .O(N__39310),
            .I(N__39301));
    Span4Mux_h I__8511 (
            .O(N__39307),
            .I(N__39301));
    InMux I__8510 (
            .O(N__39306),
            .I(N__39298));
    Odrv4 I__8509 (
            .O(N__39301),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__8508 (
            .O(N__39298),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__8507 (
            .O(N__39293),
            .I(N__39290));
    LocalMux I__8506 (
            .O(N__39290),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    InMux I__8505 (
            .O(N__39287),
            .I(N__39284));
    LocalMux I__8504 (
            .O(N__39284),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    InMux I__8503 (
            .O(N__39281),
            .I(N__39277));
    InMux I__8502 (
            .O(N__39280),
            .I(N__39274));
    LocalMux I__8501 (
            .O(N__39277),
            .I(N__39270));
    LocalMux I__8500 (
            .O(N__39274),
            .I(N__39267));
    InMux I__8499 (
            .O(N__39273),
            .I(N__39263));
    Span4Mux_h I__8498 (
            .O(N__39270),
            .I(N__39258));
    Span4Mux_h I__8497 (
            .O(N__39267),
            .I(N__39258));
    InMux I__8496 (
            .O(N__39266),
            .I(N__39255));
    LocalMux I__8495 (
            .O(N__39263),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__8494 (
            .O(N__39258),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__8493 (
            .O(N__39255),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    CascadeMux I__8492 (
            .O(N__39248),
            .I(N__39245));
    InMux I__8491 (
            .O(N__39245),
            .I(N__39242));
    LocalMux I__8490 (
            .O(N__39242),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    CascadeMux I__8489 (
            .O(N__39239),
            .I(N__39236));
    InMux I__8488 (
            .O(N__39236),
            .I(N__39231));
    InMux I__8487 (
            .O(N__39235),
            .I(N__39228));
    InMux I__8486 (
            .O(N__39234),
            .I(N__39225));
    LocalMux I__8485 (
            .O(N__39231),
            .I(N__39220));
    LocalMux I__8484 (
            .O(N__39228),
            .I(N__39220));
    LocalMux I__8483 (
            .O(N__39225),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv12 I__8482 (
            .O(N__39220),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__8481 (
            .O(N__39215),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    CascadeMux I__8480 (
            .O(N__39212),
            .I(N__39209));
    InMux I__8479 (
            .O(N__39209),
            .I(N__39202));
    InMux I__8478 (
            .O(N__39208),
            .I(N__39202));
    InMux I__8477 (
            .O(N__39207),
            .I(N__39199));
    LocalMux I__8476 (
            .O(N__39202),
            .I(N__39196));
    LocalMux I__8475 (
            .O(N__39199),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv12 I__8474 (
            .O(N__39196),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__8473 (
            .O(N__39191),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__8472 (
            .O(N__39188),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__8471 (
            .O(N__39185),
            .I(bfn_17_13_0_));
    InMux I__8470 (
            .O(N__39182),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__8469 (
            .O(N__39179),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__8468 (
            .O(N__39176),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__8467 (
            .O(N__39173),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    CascadeMux I__8466 (
            .O(N__39170),
            .I(N__39166));
    InMux I__8465 (
            .O(N__39169),
            .I(N__39160));
    InMux I__8464 (
            .O(N__39166),
            .I(N__39160));
    InMux I__8463 (
            .O(N__39165),
            .I(N__39156));
    LocalMux I__8462 (
            .O(N__39160),
            .I(N__39153));
    InMux I__8461 (
            .O(N__39159),
            .I(N__39150));
    LocalMux I__8460 (
            .O(N__39156),
            .I(N__39147));
    Span4Mux_h I__8459 (
            .O(N__39153),
            .I(N__39144));
    LocalMux I__8458 (
            .O(N__39150),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv12 I__8457 (
            .O(N__39147),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__8456 (
            .O(N__39144),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__8455 (
            .O(N__39137),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__8454 (
            .O(N__39134),
            .I(N__39130));
    InMux I__8453 (
            .O(N__39133),
            .I(N__39127));
    LocalMux I__8452 (
            .O(N__39130),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    LocalMux I__8451 (
            .O(N__39127),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__8450 (
            .O(N__39122),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__8449 (
            .O(N__39119),
            .I(N__39115));
    InMux I__8448 (
            .O(N__39118),
            .I(N__39112));
    LocalMux I__8447 (
            .O(N__39115),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__8446 (
            .O(N__39112),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__8445 (
            .O(N__39107),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__8444 (
            .O(N__39104),
            .I(N__39100));
    InMux I__8443 (
            .O(N__39103),
            .I(N__39097));
    LocalMux I__8442 (
            .O(N__39100),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__8441 (
            .O(N__39097),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__8440 (
            .O(N__39092),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__8439 (
            .O(N__39089),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__8438 (
            .O(N__39086),
            .I(bfn_17_12_0_));
    InMux I__8437 (
            .O(N__39083),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__8436 (
            .O(N__39080),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    CascadeMux I__8435 (
            .O(N__39077),
            .I(N__39073));
    InMux I__8434 (
            .O(N__39076),
            .I(N__39067));
    InMux I__8433 (
            .O(N__39073),
            .I(N__39067));
    InMux I__8432 (
            .O(N__39072),
            .I(N__39064));
    LocalMux I__8431 (
            .O(N__39067),
            .I(N__39061));
    LocalMux I__8430 (
            .O(N__39064),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__8429 (
            .O(N__39061),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__8428 (
            .O(N__39056),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__8427 (
            .O(N__39053),
            .I(N__39046));
    InMux I__8426 (
            .O(N__39052),
            .I(N__39046));
    InMux I__8425 (
            .O(N__39051),
            .I(N__39043));
    LocalMux I__8424 (
            .O(N__39046),
            .I(N__39040));
    LocalMux I__8423 (
            .O(N__39043),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__8422 (
            .O(N__39040),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__8421 (
            .O(N__39035),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__8420 (
            .O(N__39032),
            .I(N__39028));
    InMux I__8419 (
            .O(N__39031),
            .I(N__39025));
    LocalMux I__8418 (
            .O(N__39028),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__8417 (
            .O(N__39025),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__8416 (
            .O(N__39020),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__8415 (
            .O(N__39017),
            .I(N__39013));
    InMux I__8414 (
            .O(N__39016),
            .I(N__39010));
    LocalMux I__8413 (
            .O(N__39013),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__8412 (
            .O(N__39010),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__8411 (
            .O(N__39005),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__8410 (
            .O(N__39002),
            .I(N__38998));
    InMux I__8409 (
            .O(N__39001),
            .I(N__38995));
    LocalMux I__8408 (
            .O(N__38998),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__8407 (
            .O(N__38995),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__8406 (
            .O(N__38990),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__8405 (
            .O(N__38987),
            .I(N__38983));
    InMux I__8404 (
            .O(N__38986),
            .I(N__38980));
    LocalMux I__8403 (
            .O(N__38983),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__8402 (
            .O(N__38980),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__8401 (
            .O(N__38975),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__8400 (
            .O(N__38972),
            .I(N__38968));
    InMux I__8399 (
            .O(N__38971),
            .I(N__38965));
    LocalMux I__8398 (
            .O(N__38968),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__8397 (
            .O(N__38965),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__8396 (
            .O(N__38960),
            .I(bfn_17_11_0_));
    InMux I__8395 (
            .O(N__38957),
            .I(N__38953));
    InMux I__8394 (
            .O(N__38956),
            .I(N__38950));
    LocalMux I__8393 (
            .O(N__38953),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__8392 (
            .O(N__38950),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__8391 (
            .O(N__38945),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__8390 (
            .O(N__38942),
            .I(N__38938));
    InMux I__8389 (
            .O(N__38941),
            .I(N__38935));
    LocalMux I__8388 (
            .O(N__38938),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__8387 (
            .O(N__38935),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__8386 (
            .O(N__38930),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__8385 (
            .O(N__38927),
            .I(N__38923));
    InMux I__8384 (
            .O(N__38926),
            .I(N__38920));
    LocalMux I__8383 (
            .O(N__38923),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__8382 (
            .O(N__38920),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__8381 (
            .O(N__38915),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__8380 (
            .O(N__38912),
            .I(N__38907));
    InMux I__8379 (
            .O(N__38911),
            .I(N__38904));
    InMux I__8378 (
            .O(N__38910),
            .I(N__38900));
    LocalMux I__8377 (
            .O(N__38907),
            .I(N__38897));
    LocalMux I__8376 (
            .O(N__38904),
            .I(N__38894));
    InMux I__8375 (
            .O(N__38903),
            .I(N__38891));
    LocalMux I__8374 (
            .O(N__38900),
            .I(N__38888));
    Span4Mux_h I__8373 (
            .O(N__38897),
            .I(N__38885));
    Span4Mux_v I__8372 (
            .O(N__38894),
            .I(N__38880));
    LocalMux I__8371 (
            .O(N__38891),
            .I(N__38880));
    Span4Mux_h I__8370 (
            .O(N__38888),
            .I(N__38877));
    Span4Mux_v I__8369 (
            .O(N__38885),
            .I(N__38874));
    Odrv4 I__8368 (
            .O(N__38880),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv4 I__8367 (
            .O(N__38877),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv4 I__8366 (
            .O(N__38874),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__8365 (
            .O(N__38867),
            .I(N__38862));
    InMux I__8364 (
            .O(N__38866),
            .I(N__38859));
    InMux I__8363 (
            .O(N__38865),
            .I(N__38856));
    LocalMux I__8362 (
            .O(N__38862),
            .I(N__38851));
    LocalMux I__8361 (
            .O(N__38859),
            .I(N__38851));
    LocalMux I__8360 (
            .O(N__38856),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    Odrv4 I__8359 (
            .O(N__38851),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    InMux I__8358 (
            .O(N__38846),
            .I(N__38843));
    LocalMux I__8357 (
            .O(N__38843),
            .I(N__38838));
    InMux I__8356 (
            .O(N__38842),
            .I(N__38833));
    InMux I__8355 (
            .O(N__38841),
            .I(N__38833));
    Span4Mux_h I__8354 (
            .O(N__38838),
            .I(N__38830));
    LocalMux I__8353 (
            .O(N__38833),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    Odrv4 I__8352 (
            .O(N__38830),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    InMux I__8351 (
            .O(N__38825),
            .I(N__38821));
    CascadeMux I__8350 (
            .O(N__38824),
            .I(N__38818));
    LocalMux I__8349 (
            .O(N__38821),
            .I(N__38814));
    InMux I__8348 (
            .O(N__38818),
            .I(N__38809));
    InMux I__8347 (
            .O(N__38817),
            .I(N__38809));
    Span4Mux_v I__8346 (
            .O(N__38814),
            .I(N__38806));
    LocalMux I__8345 (
            .O(N__38809),
            .I(N__38801));
    Span4Mux_h I__8344 (
            .O(N__38806),
            .I(N__38801));
    Odrv4 I__8343 (
            .O(N__38801),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    InMux I__8342 (
            .O(N__38798),
            .I(N__38792));
    InMux I__8341 (
            .O(N__38797),
            .I(N__38789));
    InMux I__8340 (
            .O(N__38796),
            .I(N__38786));
    InMux I__8339 (
            .O(N__38795),
            .I(N__38783));
    LocalMux I__8338 (
            .O(N__38792),
            .I(N__38780));
    LocalMux I__8337 (
            .O(N__38789),
            .I(N__38773));
    LocalMux I__8336 (
            .O(N__38786),
            .I(N__38773));
    LocalMux I__8335 (
            .O(N__38783),
            .I(N__38773));
    Span4Mux_v I__8334 (
            .O(N__38780),
            .I(N__38770));
    Span4Mux_v I__8333 (
            .O(N__38773),
            .I(N__38767));
    Odrv4 I__8332 (
            .O(N__38770),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv4 I__8331 (
            .O(N__38767),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__8330 (
            .O(N__38762),
            .I(N__38759));
    LocalMux I__8329 (
            .O(N__38759),
            .I(N__38755));
    InMux I__8328 (
            .O(N__38758),
            .I(N__38751));
    Span4Mux_v I__8327 (
            .O(N__38755),
            .I(N__38748));
    InMux I__8326 (
            .O(N__38754),
            .I(N__38745));
    LocalMux I__8325 (
            .O(N__38751),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv4 I__8324 (
            .O(N__38748),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    LocalMux I__8323 (
            .O(N__38745),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    InMux I__8322 (
            .O(N__38738),
            .I(N__38732));
    InMux I__8321 (
            .O(N__38737),
            .I(N__38729));
    CascadeMux I__8320 (
            .O(N__38736),
            .I(N__38726));
    InMux I__8319 (
            .O(N__38735),
            .I(N__38723));
    LocalMux I__8318 (
            .O(N__38732),
            .I(N__38718));
    LocalMux I__8317 (
            .O(N__38729),
            .I(N__38718));
    InMux I__8316 (
            .O(N__38726),
            .I(N__38715));
    LocalMux I__8315 (
            .O(N__38723),
            .I(N__38712));
    Span4Mux_h I__8314 (
            .O(N__38718),
            .I(N__38709));
    LocalMux I__8313 (
            .O(N__38715),
            .I(N__38706));
    Odrv4 I__8312 (
            .O(N__38712),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__8311 (
            .O(N__38709),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__8310 (
            .O(N__38706),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__8309 (
            .O(N__38699),
            .I(N__38694));
    InMux I__8308 (
            .O(N__38698),
            .I(N__38691));
    InMux I__8307 (
            .O(N__38697),
            .I(N__38688));
    LocalMux I__8306 (
            .O(N__38694),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__8305 (
            .O(N__38691),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__8304 (
            .O(N__38688),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    CascadeMux I__8303 (
            .O(N__38681),
            .I(N__38678));
    InMux I__8302 (
            .O(N__38678),
            .I(N__38675));
    LocalMux I__8301 (
            .O(N__38675),
            .I(N__38671));
    CascadeMux I__8300 (
            .O(N__38674),
            .I(N__38667));
    Span4Mux_v I__8299 (
            .O(N__38671),
            .I(N__38664));
    InMux I__8298 (
            .O(N__38670),
            .I(N__38661));
    InMux I__8297 (
            .O(N__38667),
            .I(N__38658));
    Sp12to4 I__8296 (
            .O(N__38664),
            .I(N__38653));
    LocalMux I__8295 (
            .O(N__38661),
            .I(N__38653));
    LocalMux I__8294 (
            .O(N__38658),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv12 I__8293 (
            .O(N__38653),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__8292 (
            .O(N__38648),
            .I(N__38644));
    InMux I__8291 (
            .O(N__38647),
            .I(N__38641));
    LocalMux I__8290 (
            .O(N__38644),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__8289 (
            .O(N__38641),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__8288 (
            .O(N__38636),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    InMux I__8287 (
            .O(N__38633),
            .I(N__38629));
    InMux I__8286 (
            .O(N__38632),
            .I(N__38626));
    LocalMux I__8285 (
            .O(N__38629),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__8284 (
            .O(N__38626),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__8283 (
            .O(N__38621),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__8282 (
            .O(N__38618),
            .I(N__38614));
    InMux I__8281 (
            .O(N__38617),
            .I(N__38611));
    LocalMux I__8280 (
            .O(N__38614),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__8279 (
            .O(N__38611),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__8278 (
            .O(N__38606),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__8277 (
            .O(N__38603),
            .I(N__38600));
    LocalMux I__8276 (
            .O(N__38600),
            .I(N__38597));
    Odrv4 I__8275 (
            .O(N__38597),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ));
    InMux I__8274 (
            .O(N__38594),
            .I(N__38591));
    LocalMux I__8273 (
            .O(N__38591),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ));
    InMux I__8272 (
            .O(N__38588),
            .I(N__38585));
    LocalMux I__8271 (
            .O(N__38585),
            .I(N__38582));
    Span4Mux_h I__8270 (
            .O(N__38582),
            .I(N__38579));
    Span4Mux_v I__8269 (
            .O(N__38579),
            .I(N__38576));
    Odrv4 I__8268 (
            .O(N__38576),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt22 ));
    CascadeMux I__8267 (
            .O(N__38573),
            .I(N__38570));
    InMux I__8266 (
            .O(N__38570),
            .I(N__38567));
    LocalMux I__8265 (
            .O(N__38567),
            .I(N__38564));
    Span4Mux_v I__8264 (
            .O(N__38564),
            .I(N__38561));
    Odrv4 I__8263 (
            .O(N__38561),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ));
    InMux I__8262 (
            .O(N__38558),
            .I(N__38554));
    InMux I__8261 (
            .O(N__38557),
            .I(N__38551));
    LocalMux I__8260 (
            .O(N__38554),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__8259 (
            .O(N__38551),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    CascadeMux I__8258 (
            .O(N__38546),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_));
    InMux I__8257 (
            .O(N__38543),
            .I(N__38537));
    InMux I__8256 (
            .O(N__38542),
            .I(N__38537));
    LocalMux I__8255 (
            .O(N__38537),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ));
    InMux I__8254 (
            .O(N__38534),
            .I(N__38531));
    LocalMux I__8253 (
            .O(N__38531),
            .I(N__38528));
    Span4Mux_h I__8252 (
            .O(N__38528),
            .I(N__38525));
    Odrv4 I__8251 (
            .O(N__38525),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__8250 (
            .O(N__38522),
            .I(N__38517));
    InMux I__8249 (
            .O(N__38521),
            .I(N__38514));
    InMux I__8248 (
            .O(N__38520),
            .I(N__38511));
    InMux I__8247 (
            .O(N__38517),
            .I(N__38508));
    LocalMux I__8246 (
            .O(N__38514),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    LocalMux I__8245 (
            .O(N__38511),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    LocalMux I__8244 (
            .O(N__38508),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__8243 (
            .O(N__38501),
            .I(N__38495));
    InMux I__8242 (
            .O(N__38500),
            .I(N__38490));
    InMux I__8241 (
            .O(N__38499),
            .I(N__38490));
    InMux I__8240 (
            .O(N__38498),
            .I(N__38487));
    LocalMux I__8239 (
            .O(N__38495),
            .I(N__38482));
    LocalMux I__8238 (
            .O(N__38490),
            .I(N__38482));
    LocalMux I__8237 (
            .O(N__38487),
            .I(N__38479));
    Span4Mux_v I__8236 (
            .O(N__38482),
            .I(N__38476));
    Odrv4 I__8235 (
            .O(N__38479),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv4 I__8234 (
            .O(N__38476),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    CascadeMux I__8233 (
            .O(N__38471),
            .I(N__38468));
    InMux I__8232 (
            .O(N__38468),
            .I(N__38465));
    LocalMux I__8231 (
            .O(N__38465),
            .I(N__38462));
    Odrv4 I__8230 (
            .O(N__38462),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__8229 (
            .O(N__38459),
            .I(N__38454));
    InMux I__8228 (
            .O(N__38458),
            .I(N__38451));
    InMux I__8227 (
            .O(N__38457),
            .I(N__38448));
    InMux I__8226 (
            .O(N__38454),
            .I(N__38445));
    LocalMux I__8225 (
            .O(N__38451),
            .I(N__38439));
    LocalMux I__8224 (
            .O(N__38448),
            .I(N__38439));
    LocalMux I__8223 (
            .O(N__38445),
            .I(N__38436));
    InMux I__8222 (
            .O(N__38444),
            .I(N__38433));
    Span4Mux_v I__8221 (
            .O(N__38439),
            .I(N__38428));
    Span4Mux_v I__8220 (
            .O(N__38436),
            .I(N__38428));
    LocalMux I__8219 (
            .O(N__38433),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv4 I__8218 (
            .O(N__38428),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__8217 (
            .O(N__38423),
            .I(N__38420));
    LocalMux I__8216 (
            .O(N__38420),
            .I(N__38417));
    Odrv4 I__8215 (
            .O(N__38417),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    InMux I__8214 (
            .O(N__38414),
            .I(N__38410));
    InMux I__8213 (
            .O(N__38413),
            .I(N__38407));
    LocalMux I__8212 (
            .O(N__38410),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    LocalMux I__8211 (
            .O(N__38407),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    CascadeMux I__8210 (
            .O(N__38402),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21_cascade_));
    CascadeMux I__8209 (
            .O(N__38399),
            .I(N__38396));
    InMux I__8208 (
            .O(N__38396),
            .I(N__38390));
    InMux I__8207 (
            .O(N__38395),
            .I(N__38390));
    LocalMux I__8206 (
            .O(N__38390),
            .I(N__38387));
    Span4Mux_v I__8205 (
            .O(N__38387),
            .I(N__38384));
    Odrv4 I__8204 (
            .O(N__38384),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    CascadeMux I__8203 (
            .O(N__38381),
            .I(N__38378));
    InMux I__8202 (
            .O(N__38378),
            .I(N__38375));
    LocalMux I__8201 (
            .O(N__38375),
            .I(N__38372));
    Odrv4 I__8200 (
            .O(N__38372),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    InMux I__8199 (
            .O(N__38369),
            .I(N__38366));
    LocalMux I__8198 (
            .O(N__38366),
            .I(N__38363));
    Span4Mux_h I__8197 (
            .O(N__38363),
            .I(N__38360));
    Odrv4 I__8196 (
            .O(N__38360),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ));
    InMux I__8195 (
            .O(N__38357),
            .I(N__38353));
    InMux I__8194 (
            .O(N__38356),
            .I(N__38350));
    LocalMux I__8193 (
            .O(N__38353),
            .I(N__38347));
    LocalMux I__8192 (
            .O(N__38350),
            .I(N__38344));
    Span4Mux_h I__8191 (
            .O(N__38347),
            .I(N__38339));
    Span4Mux_h I__8190 (
            .O(N__38344),
            .I(N__38336));
    InMux I__8189 (
            .O(N__38343),
            .I(N__38331));
    InMux I__8188 (
            .O(N__38342),
            .I(N__38331));
    Span4Mux_v I__8187 (
            .O(N__38339),
            .I(N__38328));
    Odrv4 I__8186 (
            .O(N__38336),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    LocalMux I__8185 (
            .O(N__38331),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__8184 (
            .O(N__38328),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    CascadeMux I__8183 (
            .O(N__38321),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ));
    InMux I__8182 (
            .O(N__38318),
            .I(N__38315));
    LocalMux I__8181 (
            .O(N__38315),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    CascadeMux I__8180 (
            .O(N__38312),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__8179 (
            .O(N__38309),
            .I(N__38305));
    InMux I__8178 (
            .O(N__38308),
            .I(N__38302));
    LocalMux I__8177 (
            .O(N__38305),
            .I(N__38295));
    LocalMux I__8176 (
            .O(N__38302),
            .I(N__38295));
    InMux I__8175 (
            .O(N__38301),
            .I(N__38292));
    InMux I__8174 (
            .O(N__38300),
            .I(N__38289));
    Span4Mux_h I__8173 (
            .O(N__38295),
            .I(N__38286));
    LocalMux I__8172 (
            .O(N__38292),
            .I(N__38283));
    LocalMux I__8171 (
            .O(N__38289),
            .I(N__38280));
    Span4Mux_v I__8170 (
            .O(N__38286),
            .I(N__38277));
    Span4Mux_v I__8169 (
            .O(N__38283),
            .I(N__38272));
    Span4Mux_h I__8168 (
            .O(N__38280),
            .I(N__38272));
    Odrv4 I__8167 (
            .O(N__38277),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__8166 (
            .O(N__38272),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__8165 (
            .O(N__38267),
            .I(N__38259));
    InMux I__8164 (
            .O(N__38266),
            .I(N__38259));
    InMux I__8163 (
            .O(N__38265),
            .I(N__38256));
    InMux I__8162 (
            .O(N__38264),
            .I(N__38253));
    LocalMux I__8161 (
            .O(N__38259),
            .I(N__38250));
    LocalMux I__8160 (
            .O(N__38256),
            .I(N__38247));
    LocalMux I__8159 (
            .O(N__38253),
            .I(N__38244));
    Span4Mux_v I__8158 (
            .O(N__38250),
            .I(N__38241));
    Span4Mux_v I__8157 (
            .O(N__38247),
            .I(N__38236));
    Span4Mux_h I__8156 (
            .O(N__38244),
            .I(N__38236));
    Odrv4 I__8155 (
            .O(N__38241),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv4 I__8154 (
            .O(N__38236),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    CascadeMux I__8153 (
            .O(N__38231),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ));
    InMux I__8152 (
            .O(N__38228),
            .I(N__38224));
    InMux I__8151 (
            .O(N__38227),
            .I(N__38221));
    LocalMux I__8150 (
            .O(N__38224),
            .I(N__38218));
    LocalMux I__8149 (
            .O(N__38221),
            .I(N__38214));
    Span4Mux_v I__8148 (
            .O(N__38218),
            .I(N__38210));
    InMux I__8147 (
            .O(N__38217),
            .I(N__38207));
    Span4Mux_h I__8146 (
            .O(N__38214),
            .I(N__38204));
    InMux I__8145 (
            .O(N__38213),
            .I(N__38201));
    Odrv4 I__8144 (
            .O(N__38210),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__8143 (
            .O(N__38207),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    Odrv4 I__8142 (
            .O(N__38204),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__8141 (
            .O(N__38201),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__8140 (
            .O(N__38192),
            .I(N__38188));
    InMux I__8139 (
            .O(N__38191),
            .I(N__38185));
    LocalMux I__8138 (
            .O(N__38188),
            .I(N__38181));
    LocalMux I__8137 (
            .O(N__38185),
            .I(N__38178));
    InMux I__8136 (
            .O(N__38184),
            .I(N__38175));
    Span4Mux_v I__8135 (
            .O(N__38181),
            .I(N__38170));
    Span4Mux_h I__8134 (
            .O(N__38178),
            .I(N__38170));
    LocalMux I__8133 (
            .O(N__38175),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv4 I__8132 (
            .O(N__38170),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__8131 (
            .O(N__38165),
            .I(N__38162));
    LocalMux I__8130 (
            .O(N__38162),
            .I(N__38156));
    InMux I__8129 (
            .O(N__38161),
            .I(N__38153));
    InMux I__8128 (
            .O(N__38160),
            .I(N__38150));
    InMux I__8127 (
            .O(N__38159),
            .I(N__38147));
    Span4Mux_v I__8126 (
            .O(N__38156),
            .I(N__38144));
    LocalMux I__8125 (
            .O(N__38153),
            .I(N__38141));
    LocalMux I__8124 (
            .O(N__38150),
            .I(N__38138));
    LocalMux I__8123 (
            .O(N__38147),
            .I(N__38135));
    Span4Mux_v I__8122 (
            .O(N__38144),
            .I(N__38132));
    Span4Mux_h I__8121 (
            .O(N__38141),
            .I(N__38127));
    Span4Mux_h I__8120 (
            .O(N__38138),
            .I(N__38127));
    Odrv12 I__8119 (
            .O(N__38135),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    Odrv4 I__8118 (
            .O(N__38132),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    Odrv4 I__8117 (
            .O(N__38127),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__8116 (
            .O(N__38120),
            .I(N__38115));
    InMux I__8115 (
            .O(N__38119),
            .I(N__38112));
    InMux I__8114 (
            .O(N__38118),
            .I(N__38109));
    LocalMux I__8113 (
            .O(N__38115),
            .I(N__38106));
    LocalMux I__8112 (
            .O(N__38112),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    LocalMux I__8111 (
            .O(N__38109),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    Odrv4 I__8110 (
            .O(N__38106),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__8109 (
            .O(N__38099),
            .I(N__38094));
    InMux I__8108 (
            .O(N__38098),
            .I(N__38091));
    InMux I__8107 (
            .O(N__38097),
            .I(N__38088));
    LocalMux I__8106 (
            .O(N__38094),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    LocalMux I__8105 (
            .O(N__38091),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    LocalMux I__8104 (
            .O(N__38088),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    InMux I__8103 (
            .O(N__38081),
            .I(N__38076));
    InMux I__8102 (
            .O(N__38080),
            .I(N__38073));
    InMux I__8101 (
            .O(N__38079),
            .I(N__38070));
    LocalMux I__8100 (
            .O(N__38076),
            .I(N__38067));
    LocalMux I__8099 (
            .O(N__38073),
            .I(\phase_controller_inst1.tr_time_passed ));
    LocalMux I__8098 (
            .O(N__38070),
            .I(\phase_controller_inst1.tr_time_passed ));
    Odrv4 I__8097 (
            .O(N__38067),
            .I(\phase_controller_inst1.tr_time_passed ));
    CascadeMux I__8096 (
            .O(N__38060),
            .I(N__38057));
    InMux I__8095 (
            .O(N__38057),
            .I(N__38050));
    InMux I__8094 (
            .O(N__38056),
            .I(N__38050));
    InMux I__8093 (
            .O(N__38055),
            .I(N__38047));
    LocalMux I__8092 (
            .O(N__38050),
            .I(N__38043));
    LocalMux I__8091 (
            .O(N__38047),
            .I(N__38040));
    InMux I__8090 (
            .O(N__38046),
            .I(N__38037));
    Span4Mux_v I__8089 (
            .O(N__38043),
            .I(N__38034));
    Span4Mux_h I__8088 (
            .O(N__38040),
            .I(N__38031));
    LocalMux I__8087 (
            .O(N__38037),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    Odrv4 I__8086 (
            .O(N__38034),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    Odrv4 I__8085 (
            .O(N__38031),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__8084 (
            .O(N__38024),
            .I(N__38021));
    LocalMux I__8083 (
            .O(N__38021),
            .I(N__38017));
    InMux I__8082 (
            .O(N__38020),
            .I(N__38014));
    Span4Mux_v I__8081 (
            .O(N__38017),
            .I(N__38011));
    LocalMux I__8080 (
            .O(N__38014),
            .I(N__38008));
    Odrv4 I__8079 (
            .O(N__38011),
            .I(\phase_controller_inst1.time_passed_RNI7NN7 ));
    Odrv4 I__8078 (
            .O(N__38008),
            .I(\phase_controller_inst1.time_passed_RNI7NN7 ));
    InMux I__8077 (
            .O(N__38003),
            .I(N__37987));
    InMux I__8076 (
            .O(N__38002),
            .I(N__37984));
    InMux I__8075 (
            .O(N__38001),
            .I(N__37981));
    CascadeMux I__8074 (
            .O(N__38000),
            .I(N__37972));
    CascadeMux I__8073 (
            .O(N__37999),
            .I(N__37968));
    CascadeMux I__8072 (
            .O(N__37998),
            .I(N__37964));
    CascadeMux I__8071 (
            .O(N__37997),
            .I(N__37960));
    CascadeMux I__8070 (
            .O(N__37996),
            .I(N__37956));
    CascadeMux I__8069 (
            .O(N__37995),
            .I(N__37952));
    CascadeMux I__8068 (
            .O(N__37994),
            .I(N__37948));
    CascadeMux I__8067 (
            .O(N__37993),
            .I(N__37944));
    CascadeMux I__8066 (
            .O(N__37992),
            .I(N__37940));
    CascadeMux I__8065 (
            .O(N__37991),
            .I(N__37936));
    CascadeMux I__8064 (
            .O(N__37990),
            .I(N__37932));
    LocalMux I__8063 (
            .O(N__37987),
            .I(N__37921));
    LocalMux I__8062 (
            .O(N__37984),
            .I(N__37921));
    LocalMux I__8061 (
            .O(N__37981),
            .I(N__37921));
    InMux I__8060 (
            .O(N__37980),
            .I(N__37918));
    InMux I__8059 (
            .O(N__37979),
            .I(N__37914));
    InMux I__8058 (
            .O(N__37978),
            .I(N__37909));
    InMux I__8057 (
            .O(N__37977),
            .I(N__37909));
    InMux I__8056 (
            .O(N__37976),
            .I(N__37906));
    InMux I__8055 (
            .O(N__37975),
            .I(N__37894));
    InMux I__8054 (
            .O(N__37972),
            .I(N__37879));
    InMux I__8053 (
            .O(N__37971),
            .I(N__37879));
    InMux I__8052 (
            .O(N__37968),
            .I(N__37879));
    InMux I__8051 (
            .O(N__37967),
            .I(N__37879));
    InMux I__8050 (
            .O(N__37964),
            .I(N__37879));
    InMux I__8049 (
            .O(N__37963),
            .I(N__37879));
    InMux I__8048 (
            .O(N__37960),
            .I(N__37879));
    InMux I__8047 (
            .O(N__37959),
            .I(N__37864));
    InMux I__8046 (
            .O(N__37956),
            .I(N__37864));
    InMux I__8045 (
            .O(N__37955),
            .I(N__37864));
    InMux I__8044 (
            .O(N__37952),
            .I(N__37864));
    InMux I__8043 (
            .O(N__37951),
            .I(N__37864));
    InMux I__8042 (
            .O(N__37948),
            .I(N__37864));
    InMux I__8041 (
            .O(N__37947),
            .I(N__37864));
    InMux I__8040 (
            .O(N__37944),
            .I(N__37847));
    InMux I__8039 (
            .O(N__37943),
            .I(N__37847));
    InMux I__8038 (
            .O(N__37940),
            .I(N__37847));
    InMux I__8037 (
            .O(N__37939),
            .I(N__37847));
    InMux I__8036 (
            .O(N__37936),
            .I(N__37847));
    InMux I__8035 (
            .O(N__37935),
            .I(N__37847));
    InMux I__8034 (
            .O(N__37932),
            .I(N__37847));
    InMux I__8033 (
            .O(N__37931),
            .I(N__37847));
    InMux I__8032 (
            .O(N__37930),
            .I(N__37840));
    InMux I__8031 (
            .O(N__37929),
            .I(N__37835));
    InMux I__8030 (
            .O(N__37928),
            .I(N__37835));
    Span4Mux_s2_v I__8029 (
            .O(N__37921),
            .I(N__37830));
    LocalMux I__8028 (
            .O(N__37918),
            .I(N__37830));
    CascadeMux I__8027 (
            .O(N__37917),
            .I(N__37819));
    LocalMux I__8026 (
            .O(N__37914),
            .I(N__37815));
    LocalMux I__8025 (
            .O(N__37909),
            .I(N__37810));
    LocalMux I__8024 (
            .O(N__37906),
            .I(N__37810));
    InMux I__8023 (
            .O(N__37905),
            .I(N__37807));
    InMux I__8022 (
            .O(N__37904),
            .I(N__37804));
    InMux I__8021 (
            .O(N__37903),
            .I(N__37797));
    InMux I__8020 (
            .O(N__37902),
            .I(N__37797));
    InMux I__8019 (
            .O(N__37901),
            .I(N__37797));
    InMux I__8018 (
            .O(N__37900),
            .I(N__37788));
    InMux I__8017 (
            .O(N__37899),
            .I(N__37788));
    InMux I__8016 (
            .O(N__37898),
            .I(N__37788));
    InMux I__8015 (
            .O(N__37897),
            .I(N__37788));
    LocalMux I__8014 (
            .O(N__37894),
            .I(N__37785));
    LocalMux I__8013 (
            .O(N__37879),
            .I(N__37782));
    LocalMux I__8012 (
            .O(N__37864),
            .I(N__37777));
    LocalMux I__8011 (
            .O(N__37847),
            .I(N__37777));
    CascadeMux I__8010 (
            .O(N__37846),
            .I(N__37774));
    CascadeMux I__8009 (
            .O(N__37845),
            .I(N__37770));
    CascadeMux I__8008 (
            .O(N__37844),
            .I(N__37766));
    CascadeMux I__8007 (
            .O(N__37843),
            .I(N__37762));
    LocalMux I__8006 (
            .O(N__37840),
            .I(N__37756));
    LocalMux I__8005 (
            .O(N__37835),
            .I(N__37753));
    Span4Mux_v I__8004 (
            .O(N__37830),
            .I(N__37750));
    InMux I__8003 (
            .O(N__37829),
            .I(N__37743));
    InMux I__8002 (
            .O(N__37828),
            .I(N__37743));
    InMux I__8001 (
            .O(N__37827),
            .I(N__37743));
    InMux I__8000 (
            .O(N__37826),
            .I(N__37734));
    InMux I__7999 (
            .O(N__37825),
            .I(N__37734));
    InMux I__7998 (
            .O(N__37824),
            .I(N__37734));
    InMux I__7997 (
            .O(N__37823),
            .I(N__37734));
    InMux I__7996 (
            .O(N__37822),
            .I(N__37727));
    InMux I__7995 (
            .O(N__37819),
            .I(N__37727));
    InMux I__7994 (
            .O(N__37818),
            .I(N__37727));
    Span4Mux_v I__7993 (
            .O(N__37815),
            .I(N__37720));
    Span4Mux_v I__7992 (
            .O(N__37810),
            .I(N__37720));
    LocalMux I__7991 (
            .O(N__37807),
            .I(N__37720));
    LocalMux I__7990 (
            .O(N__37804),
            .I(N__37711));
    LocalMux I__7989 (
            .O(N__37797),
            .I(N__37711));
    LocalMux I__7988 (
            .O(N__37788),
            .I(N__37711));
    Span12Mux_s2_v I__7987 (
            .O(N__37785),
            .I(N__37711));
    Span4Mux_v I__7986 (
            .O(N__37782),
            .I(N__37706));
    Span4Mux_v I__7985 (
            .O(N__37777),
            .I(N__37706));
    InMux I__7984 (
            .O(N__37774),
            .I(N__37689));
    InMux I__7983 (
            .O(N__37773),
            .I(N__37689));
    InMux I__7982 (
            .O(N__37770),
            .I(N__37689));
    InMux I__7981 (
            .O(N__37769),
            .I(N__37689));
    InMux I__7980 (
            .O(N__37766),
            .I(N__37689));
    InMux I__7979 (
            .O(N__37765),
            .I(N__37689));
    InMux I__7978 (
            .O(N__37762),
            .I(N__37689));
    InMux I__7977 (
            .O(N__37761),
            .I(N__37689));
    InMux I__7976 (
            .O(N__37760),
            .I(N__37684));
    InMux I__7975 (
            .O(N__37759),
            .I(N__37684));
    Span4Mux_s1_h I__7974 (
            .O(N__37756),
            .I(N__37679));
    Span4Mux_v I__7973 (
            .O(N__37753),
            .I(N__37679));
    Sp12to4 I__7972 (
            .O(N__37750),
            .I(N__37670));
    LocalMux I__7971 (
            .O(N__37743),
            .I(N__37670));
    LocalMux I__7970 (
            .O(N__37734),
            .I(N__37670));
    LocalMux I__7969 (
            .O(N__37727),
            .I(N__37670));
    Sp12to4 I__7968 (
            .O(N__37720),
            .I(N__37667));
    Span12Mux_v I__7967 (
            .O(N__37711),
            .I(N__37660));
    Sp12to4 I__7966 (
            .O(N__37706),
            .I(N__37660));
    LocalMux I__7965 (
            .O(N__37689),
            .I(N__37660));
    LocalMux I__7964 (
            .O(N__37684),
            .I(N__37657));
    Span4Mux_h I__7963 (
            .O(N__37679),
            .I(N__37654));
    Span12Mux_s5_h I__7962 (
            .O(N__37670),
            .I(N__37651));
    Span12Mux_v I__7961 (
            .O(N__37667),
            .I(N__37644));
    Span12Mux_h I__7960 (
            .O(N__37660),
            .I(N__37644));
    Span12Mux_v I__7959 (
            .O(N__37657),
            .I(N__37644));
    Odrv4 I__7958 (
            .O(N__37654),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__7957 (
            .O(N__37651),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__7956 (
            .O(N__37644),
            .I(CONSTANT_ONE_NET));
    InMux I__7955 (
            .O(N__37637),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__7954 (
            .O(N__37634),
            .I(N__37628));
    CascadeMux I__7953 (
            .O(N__37633),
            .I(N__37625));
    InMux I__7952 (
            .O(N__37632),
            .I(N__37616));
    InMux I__7951 (
            .O(N__37631),
            .I(N__37616));
    LocalMux I__7950 (
            .O(N__37628),
            .I(N__37613));
    InMux I__7949 (
            .O(N__37625),
            .I(N__37610));
    InMux I__7948 (
            .O(N__37624),
            .I(N__37607));
    InMux I__7947 (
            .O(N__37623),
            .I(N__37602));
    InMux I__7946 (
            .O(N__37622),
            .I(N__37602));
    CascadeMux I__7945 (
            .O(N__37621),
            .I(N__37595));
    LocalMux I__7944 (
            .O(N__37616),
            .I(N__37590));
    Span4Mux_v I__7943 (
            .O(N__37613),
            .I(N__37586));
    LocalMux I__7942 (
            .O(N__37610),
            .I(N__37583));
    LocalMux I__7941 (
            .O(N__37607),
            .I(N__37578));
    LocalMux I__7940 (
            .O(N__37602),
            .I(N__37578));
    InMux I__7939 (
            .O(N__37601),
            .I(N__37563));
    InMux I__7938 (
            .O(N__37600),
            .I(N__37563));
    InMux I__7937 (
            .O(N__37599),
            .I(N__37563));
    InMux I__7936 (
            .O(N__37598),
            .I(N__37563));
    InMux I__7935 (
            .O(N__37595),
            .I(N__37563));
    InMux I__7934 (
            .O(N__37594),
            .I(N__37563));
    InMux I__7933 (
            .O(N__37593),
            .I(N__37563));
    Span4Mux_h I__7932 (
            .O(N__37590),
            .I(N__37560));
    InMux I__7931 (
            .O(N__37589),
            .I(N__37557));
    Span4Mux_h I__7930 (
            .O(N__37586),
            .I(N__37552));
    Span4Mux_v I__7929 (
            .O(N__37583),
            .I(N__37552));
    Span4Mux_v I__7928 (
            .O(N__37578),
            .I(N__37547));
    LocalMux I__7927 (
            .O(N__37563),
            .I(N__37547));
    Span4Mux_h I__7926 (
            .O(N__37560),
            .I(N__37544));
    LocalMux I__7925 (
            .O(N__37557),
            .I(N__37541));
    Odrv4 I__7924 (
            .O(N__37552),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__7923 (
            .O(N__37547),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__7922 (
            .O(N__37544),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv12 I__7921 (
            .O(N__37541),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__7920 (
            .O(N__37532),
            .I(N__37529));
    LocalMux I__7919 (
            .O(N__37529),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    CascadeMux I__7918 (
            .O(N__37526),
            .I(N__37523));
    InMux I__7917 (
            .O(N__37523),
            .I(N__37520));
    LocalMux I__7916 (
            .O(N__37520),
            .I(N__37517));
    Span4Mux_v I__7915 (
            .O(N__37517),
            .I(N__37514));
    Odrv4 I__7914 (
            .O(N__37514),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ));
    InMux I__7913 (
            .O(N__37511),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ));
    InMux I__7912 (
            .O(N__37508),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ));
    CascadeMux I__7911 (
            .O(N__37505),
            .I(N__37502));
    InMux I__7910 (
            .O(N__37502),
            .I(N__37498));
    InMux I__7909 (
            .O(N__37501),
            .I(N__37495));
    LocalMux I__7908 (
            .O(N__37498),
            .I(N__37492));
    LocalMux I__7907 (
            .O(N__37495),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    Odrv12 I__7906 (
            .O(N__37492),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    CascadeMux I__7905 (
            .O(N__37487),
            .I(N__37484));
    InMux I__7904 (
            .O(N__37484),
            .I(N__37481));
    LocalMux I__7903 (
            .O(N__37481),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    CascadeMux I__7902 (
            .O(N__37478),
            .I(N__37475));
    InMux I__7901 (
            .O(N__37475),
            .I(N__37472));
    LocalMux I__7900 (
            .O(N__37472),
            .I(N__37469));
    Odrv4 I__7899 (
            .O(N__37469),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__7898 (
            .O(N__37466),
            .I(N__37463));
    InMux I__7897 (
            .O(N__37463),
            .I(N__37460));
    LocalMux I__7896 (
            .O(N__37460),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__7895 (
            .O(N__37457),
            .I(N__37454));
    LocalMux I__7894 (
            .O(N__37454),
            .I(N__37451));
    Odrv4 I__7893 (
            .O(N__37451),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ));
    CascadeMux I__7892 (
            .O(N__37448),
            .I(N__37445));
    InMux I__7891 (
            .O(N__37445),
            .I(N__37442));
    LocalMux I__7890 (
            .O(N__37442),
            .I(N__37439));
    Span4Mux_v I__7889 (
            .O(N__37439),
            .I(N__37436));
    Odrv4 I__7888 (
            .O(N__37436),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt20 ));
    InMux I__7887 (
            .O(N__37433),
            .I(N__37430));
    LocalMux I__7886 (
            .O(N__37430),
            .I(N__37427));
    Odrv12 I__7885 (
            .O(N__37427),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__7884 (
            .O(N__37424),
            .I(N__37421));
    InMux I__7883 (
            .O(N__37421),
            .I(N__37418));
    LocalMux I__7882 (
            .O(N__37418),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    CascadeMux I__7881 (
            .O(N__37415),
            .I(N__37412));
    InMux I__7880 (
            .O(N__37412),
            .I(N__37409));
    LocalMux I__7879 (
            .O(N__37409),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__7878 (
            .O(N__37406),
            .I(N__37403));
    LocalMux I__7877 (
            .O(N__37403),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__7876 (
            .O(N__37400),
            .I(N__37397));
    LocalMux I__7875 (
            .O(N__37397),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    CascadeMux I__7874 (
            .O(N__37394),
            .I(N__37391));
    InMux I__7873 (
            .O(N__37391),
            .I(N__37388));
    LocalMux I__7872 (
            .O(N__37388),
            .I(N__37385));
    Odrv4 I__7871 (
            .O(N__37385),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    InMux I__7870 (
            .O(N__37382),
            .I(N__37379));
    LocalMux I__7869 (
            .O(N__37379),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__7868 (
            .O(N__37376),
            .I(N__37373));
    LocalMux I__7867 (
            .O(N__37373),
            .I(N__37370));
    Odrv12 I__7866 (
            .O(N__37370),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__7865 (
            .O(N__37367),
            .I(N__37364));
    InMux I__7864 (
            .O(N__37364),
            .I(N__37361));
    LocalMux I__7863 (
            .O(N__37361),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__7862 (
            .O(N__37358),
            .I(N__37355));
    LocalMux I__7861 (
            .O(N__37355),
            .I(N__37352));
    Odrv4 I__7860 (
            .O(N__37352),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__7859 (
            .O(N__37349),
            .I(N__37346));
    InMux I__7858 (
            .O(N__37346),
            .I(N__37343));
    LocalMux I__7857 (
            .O(N__37343),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    CascadeMux I__7856 (
            .O(N__37340),
            .I(N__37337));
    InMux I__7855 (
            .O(N__37337),
            .I(N__37334));
    LocalMux I__7854 (
            .O(N__37334),
            .I(N__37331));
    Odrv4 I__7853 (
            .O(N__37331),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    InMux I__7852 (
            .O(N__37328),
            .I(N__37325));
    LocalMux I__7851 (
            .O(N__37325),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    InMux I__7850 (
            .O(N__37322),
            .I(N__37316));
    InMux I__7849 (
            .O(N__37321),
            .I(N__37316));
    LocalMux I__7848 (
            .O(N__37316),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    InMux I__7847 (
            .O(N__37313),
            .I(N__37310));
    LocalMux I__7846 (
            .O(N__37310),
            .I(N__37306));
    InMux I__7845 (
            .O(N__37309),
            .I(N__37302));
    Span4Mux_v I__7844 (
            .O(N__37306),
            .I(N__37299));
    InMux I__7843 (
            .O(N__37305),
            .I(N__37296));
    LocalMux I__7842 (
            .O(N__37302),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__7841 (
            .O(N__37299),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    LocalMux I__7840 (
            .O(N__37296),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__7839 (
            .O(N__37289),
            .I(N__37286));
    LocalMux I__7838 (
            .O(N__37286),
            .I(N__37283));
    Span4Mux_v I__7837 (
            .O(N__37283),
            .I(N__37277));
    InMux I__7836 (
            .O(N__37282),
            .I(N__37274));
    InMux I__7835 (
            .O(N__37281),
            .I(N__37269));
    InMux I__7834 (
            .O(N__37280),
            .I(N__37269));
    Odrv4 I__7833 (
            .O(N__37277),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__7832 (
            .O(N__37274),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    LocalMux I__7831 (
            .O(N__37269),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    CascadeMux I__7830 (
            .O(N__37262),
            .I(N__37257));
    InMux I__7829 (
            .O(N__37261),
            .I(N__37254));
    InMux I__7828 (
            .O(N__37260),
            .I(N__37251));
    InMux I__7827 (
            .O(N__37257),
            .I(N__37248));
    LocalMux I__7826 (
            .O(N__37254),
            .I(N__37244));
    LocalMux I__7825 (
            .O(N__37251),
            .I(N__37241));
    LocalMux I__7824 (
            .O(N__37248),
            .I(N__37238));
    InMux I__7823 (
            .O(N__37247),
            .I(N__37235));
    Span4Mux_v I__7822 (
            .O(N__37244),
            .I(N__37230));
    Span4Mux_h I__7821 (
            .O(N__37241),
            .I(N__37230));
    Span4Mux_h I__7820 (
            .O(N__37238),
            .I(N__37227));
    LocalMux I__7819 (
            .O(N__37235),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv4 I__7818 (
            .O(N__37230),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv4 I__7817 (
            .O(N__37227),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__7816 (
            .O(N__37220),
            .I(N__37217));
    LocalMux I__7815 (
            .O(N__37217),
            .I(N__37213));
    InMux I__7814 (
            .O(N__37216),
            .I(N__37209));
    Span4Mux_h I__7813 (
            .O(N__37213),
            .I(N__37206));
    InMux I__7812 (
            .O(N__37212),
            .I(N__37203));
    LocalMux I__7811 (
            .O(N__37209),
            .I(N__37198));
    Span4Mux_h I__7810 (
            .O(N__37206),
            .I(N__37198));
    LocalMux I__7809 (
            .O(N__37203),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    Odrv4 I__7808 (
            .O(N__37198),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    CascadeMux I__7807 (
            .O(N__37193),
            .I(N__37190));
    InMux I__7806 (
            .O(N__37190),
            .I(N__37187));
    LocalMux I__7805 (
            .O(N__37187),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    InMux I__7804 (
            .O(N__37184),
            .I(N__37181));
    LocalMux I__7803 (
            .O(N__37181),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__7802 (
            .O(N__37178),
            .I(N__37175));
    LocalMux I__7801 (
            .O(N__37175),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__7800 (
            .O(N__37172),
            .I(N__37169));
    InMux I__7799 (
            .O(N__37169),
            .I(N__37166));
    LocalMux I__7798 (
            .O(N__37166),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__7797 (
            .O(N__37163),
            .I(N__37160));
    LocalMux I__7796 (
            .O(N__37160),
            .I(N__37157));
    Span4Mux_v I__7795 (
            .O(N__37157),
            .I(N__37154));
    Odrv4 I__7794 (
            .O(N__37154),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__7793 (
            .O(N__37151),
            .I(N__37148));
    InMux I__7792 (
            .O(N__37148),
            .I(N__37145));
    LocalMux I__7791 (
            .O(N__37145),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    CascadeMux I__7790 (
            .O(N__37142),
            .I(N__37139));
    InMux I__7789 (
            .O(N__37139),
            .I(N__37136));
    LocalMux I__7788 (
            .O(N__37136),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    InMux I__7787 (
            .O(N__37133),
            .I(N__37130));
    LocalMux I__7786 (
            .O(N__37130),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__7785 (
            .O(N__37127),
            .I(N__37124));
    LocalMux I__7784 (
            .O(N__37124),
            .I(N__37121));
    Span4Mux_v I__7783 (
            .O(N__37121),
            .I(N__37118));
    Odrv4 I__7782 (
            .O(N__37118),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__7781 (
            .O(N__37115),
            .I(N__37112));
    InMux I__7780 (
            .O(N__37112),
            .I(N__37109));
    LocalMux I__7779 (
            .O(N__37109),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__7778 (
            .O(N__37106),
            .I(N__37103));
    InMux I__7777 (
            .O(N__37103),
            .I(N__37100));
    LocalMux I__7776 (
            .O(N__37100),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    InMux I__7775 (
            .O(N__37097),
            .I(N__37093));
    InMux I__7774 (
            .O(N__37096),
            .I(N__37090));
    LocalMux I__7773 (
            .O(N__37093),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__7772 (
            .O(N__37090),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    CascadeMux I__7771 (
            .O(N__37085),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_));
    InMux I__7770 (
            .O(N__37082),
            .I(N__37079));
    LocalMux I__7769 (
            .O(N__37079),
            .I(N__37075));
    InMux I__7768 (
            .O(N__37078),
            .I(N__37072));
    Odrv4 I__7767 (
            .O(N__37075),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__7766 (
            .O(N__37072),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    CascadeMux I__7765 (
            .O(N__37067),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_));
    InMux I__7764 (
            .O(N__37064),
            .I(N__37061));
    LocalMux I__7763 (
            .O(N__37061),
            .I(N__37055));
    InMux I__7762 (
            .O(N__37060),
            .I(N__37048));
    InMux I__7761 (
            .O(N__37059),
            .I(N__37048));
    InMux I__7760 (
            .O(N__37058),
            .I(N__37048));
    Span4Mux_h I__7759 (
            .O(N__37055),
            .I(N__37043));
    LocalMux I__7758 (
            .O(N__37048),
            .I(N__37043));
    Odrv4 I__7757 (
            .O(N__37043),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__7756 (
            .O(N__37040),
            .I(N__37037));
    LocalMux I__7755 (
            .O(N__37037),
            .I(N__37034));
    Span4Mux_h I__7754 (
            .O(N__37034),
            .I(N__37028));
    InMux I__7753 (
            .O(N__37033),
            .I(N__37021));
    InMux I__7752 (
            .O(N__37032),
            .I(N__37021));
    InMux I__7751 (
            .O(N__37031),
            .I(N__37021));
    Odrv4 I__7750 (
            .O(N__37028),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__7749 (
            .O(N__37021),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__7748 (
            .O(N__37016),
            .I(N__37010));
    InMux I__7747 (
            .O(N__37015),
            .I(N__37010));
    LocalMux I__7746 (
            .O(N__37010),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    InMux I__7745 (
            .O(N__37007),
            .I(N__37004));
    LocalMux I__7744 (
            .O(N__37004),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__7743 (
            .O(N__37001),
            .I(N__36998));
    InMux I__7742 (
            .O(N__36998),
            .I(N__36995));
    LocalMux I__7741 (
            .O(N__36995),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    InMux I__7740 (
            .O(N__36992),
            .I(N__36989));
    LocalMux I__7739 (
            .O(N__36989),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__7738 (
            .O(N__36986),
            .I(N__36983));
    InMux I__7737 (
            .O(N__36983),
            .I(N__36980));
    LocalMux I__7736 (
            .O(N__36980),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt22 ));
    InMux I__7735 (
            .O(N__36977),
            .I(N__36971));
    InMux I__7734 (
            .O(N__36976),
            .I(N__36971));
    LocalMux I__7733 (
            .O(N__36971),
            .I(N__36967));
    InMux I__7732 (
            .O(N__36970),
            .I(N__36964));
    Span4Mux_h I__7731 (
            .O(N__36967),
            .I(N__36961));
    LocalMux I__7730 (
            .O(N__36964),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__7729 (
            .O(N__36961),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    CascadeMux I__7728 (
            .O(N__36956),
            .I(N__36953));
    InMux I__7727 (
            .O(N__36953),
            .I(N__36947));
    InMux I__7726 (
            .O(N__36952),
            .I(N__36947));
    LocalMux I__7725 (
            .O(N__36947),
            .I(N__36943));
    InMux I__7724 (
            .O(N__36946),
            .I(N__36940));
    Span4Mux_v I__7723 (
            .O(N__36943),
            .I(N__36937));
    LocalMux I__7722 (
            .O(N__36940),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__7721 (
            .O(N__36937),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__7720 (
            .O(N__36932),
            .I(N__36929));
    LocalMux I__7719 (
            .O(N__36929),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ));
    InMux I__7718 (
            .O(N__36926),
            .I(N__36920));
    InMux I__7717 (
            .O(N__36925),
            .I(N__36920));
    LocalMux I__7716 (
            .O(N__36920),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ));
    CascadeMux I__7715 (
            .O(N__36917),
            .I(N__36914));
    InMux I__7714 (
            .O(N__36914),
            .I(N__36908));
    InMux I__7713 (
            .O(N__36913),
            .I(N__36908));
    LocalMux I__7712 (
            .O(N__36908),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ));
    CascadeMux I__7711 (
            .O(N__36905),
            .I(N__36902));
    InMux I__7710 (
            .O(N__36902),
            .I(N__36899));
    LocalMux I__7709 (
            .O(N__36899),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    InMux I__7708 (
            .O(N__36896),
            .I(N__36893));
    LocalMux I__7707 (
            .O(N__36893),
            .I(N__36890));
    Span4Mux_h I__7706 (
            .O(N__36890),
            .I(N__36885));
    InMux I__7705 (
            .O(N__36889),
            .I(N__36880));
    InMux I__7704 (
            .O(N__36888),
            .I(N__36880));
    Odrv4 I__7703 (
            .O(N__36885),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    LocalMux I__7702 (
            .O(N__36880),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    InMux I__7701 (
            .O(N__36875),
            .I(N__36872));
    LocalMux I__7700 (
            .O(N__36872),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    InMux I__7699 (
            .O(N__36869),
            .I(N__36866));
    LocalMux I__7698 (
            .O(N__36866),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    InMux I__7697 (
            .O(N__36863),
            .I(N__36859));
    InMux I__7696 (
            .O(N__36862),
            .I(N__36856));
    LocalMux I__7695 (
            .O(N__36859),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    LocalMux I__7694 (
            .O(N__36856),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__7693 (
            .O(N__36851),
            .I(N__36848));
    InMux I__7692 (
            .O(N__36848),
            .I(N__36845));
    LocalMux I__7691 (
            .O(N__36845),
            .I(N__36842));
    Span4Mux_h I__7690 (
            .O(N__36842),
            .I(N__36839));
    Odrv4 I__7689 (
            .O(N__36839),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt20 ));
    InMux I__7688 (
            .O(N__36836),
            .I(N__36830));
    InMux I__7687 (
            .O(N__36835),
            .I(N__36830));
    LocalMux I__7686 (
            .O(N__36830),
            .I(N__36826));
    InMux I__7685 (
            .O(N__36829),
            .I(N__36823));
    Span4Mux_h I__7684 (
            .O(N__36826),
            .I(N__36820));
    LocalMux I__7683 (
            .O(N__36823),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__7682 (
            .O(N__36820),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    CascadeMux I__7681 (
            .O(N__36815),
            .I(N__36811));
    CascadeMux I__7680 (
            .O(N__36814),
            .I(N__36808));
    InMux I__7679 (
            .O(N__36811),
            .I(N__36805));
    InMux I__7678 (
            .O(N__36808),
            .I(N__36802));
    LocalMux I__7677 (
            .O(N__36805),
            .I(N__36796));
    LocalMux I__7676 (
            .O(N__36802),
            .I(N__36796));
    InMux I__7675 (
            .O(N__36801),
            .I(N__36793));
    Span4Mux_v I__7674 (
            .O(N__36796),
            .I(N__36790));
    LocalMux I__7673 (
            .O(N__36793),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__7672 (
            .O(N__36790),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__7671 (
            .O(N__36785),
            .I(N__36781));
    InMux I__7670 (
            .O(N__36784),
            .I(N__36778));
    LocalMux I__7669 (
            .O(N__36781),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    LocalMux I__7668 (
            .O(N__36778),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    InMux I__7667 (
            .O(N__36773),
            .I(N__36770));
    LocalMux I__7666 (
            .O(N__36770),
            .I(N__36767));
    Odrv4 I__7665 (
            .O(N__36767),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ));
    InMux I__7664 (
            .O(N__36764),
            .I(bfn_15_21_0_));
    InMux I__7663 (
            .O(N__36761),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__7662 (
            .O(N__36758),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__7661 (
            .O(N__36755),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__7660 (
            .O(N__36752),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    IoInMux I__7659 (
            .O(N__36749),
            .I(N__36746));
    LocalMux I__7658 (
            .O(N__36746),
            .I(N__36743));
    Span4Mux_s3_v I__7657 (
            .O(N__36743),
            .I(N__36740));
    Span4Mux_v I__7656 (
            .O(N__36740),
            .I(N__36736));
    InMux I__7655 (
            .O(N__36739),
            .I(N__36733));
    Odrv4 I__7654 (
            .O(N__36736),
            .I(T12_c));
    LocalMux I__7653 (
            .O(N__36733),
            .I(T12_c));
    IoInMux I__7652 (
            .O(N__36728),
            .I(N__36725));
    LocalMux I__7651 (
            .O(N__36725),
            .I(N__36722));
    Span4Mux_s3_v I__7650 (
            .O(N__36722),
            .I(N__36718));
    InMux I__7649 (
            .O(N__36721),
            .I(N__36715));
    Odrv4 I__7648 (
            .O(N__36718),
            .I(T45_c));
    LocalMux I__7647 (
            .O(N__36715),
            .I(T45_c));
    InMux I__7646 (
            .O(N__36710),
            .I(N__36704));
    InMux I__7645 (
            .O(N__36709),
            .I(N__36704));
    LocalMux I__7644 (
            .O(N__36704),
            .I(N__36700));
    InMux I__7643 (
            .O(N__36703),
            .I(N__36697));
    Span4Mux_h I__7642 (
            .O(N__36700),
            .I(N__36690));
    LocalMux I__7641 (
            .O(N__36697),
            .I(N__36687));
    InMux I__7640 (
            .O(N__36696),
            .I(N__36684));
    InMux I__7639 (
            .O(N__36695),
            .I(N__36679));
    InMux I__7638 (
            .O(N__36694),
            .I(N__36679));
    InMux I__7637 (
            .O(N__36693),
            .I(N__36675));
    Span4Mux_v I__7636 (
            .O(N__36690),
            .I(N__36672));
    Span4Mux_v I__7635 (
            .O(N__36687),
            .I(N__36669));
    LocalMux I__7634 (
            .O(N__36684),
            .I(N__36664));
    LocalMux I__7633 (
            .O(N__36679),
            .I(N__36664));
    InMux I__7632 (
            .O(N__36678),
            .I(N__36661));
    LocalMux I__7631 (
            .O(N__36675),
            .I(state_3));
    Odrv4 I__7630 (
            .O(N__36672),
            .I(state_3));
    Odrv4 I__7629 (
            .O(N__36669),
            .I(state_3));
    Odrv12 I__7628 (
            .O(N__36664),
            .I(state_3));
    LocalMux I__7627 (
            .O(N__36661),
            .I(state_3));
    InMux I__7626 (
            .O(N__36650),
            .I(N__36646));
    InMux I__7625 (
            .O(N__36649),
            .I(N__36643));
    LocalMux I__7624 (
            .O(N__36646),
            .I(N__36640));
    LocalMux I__7623 (
            .O(N__36643),
            .I(N__36637));
    Span4Mux_h I__7622 (
            .O(N__36640),
            .I(N__36631));
    Span4Mux_h I__7621 (
            .O(N__36637),
            .I(N__36628));
    InMux I__7620 (
            .O(N__36636),
            .I(N__36625));
    InMux I__7619 (
            .O(N__36635),
            .I(N__36622));
    InMux I__7618 (
            .O(N__36634),
            .I(N__36619));
    Odrv4 I__7617 (
            .O(N__36631),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__7616 (
            .O(N__36628),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__7615 (
            .O(N__36625),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__7614 (
            .O(N__36622),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__7613 (
            .O(N__36619),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    IoInMux I__7612 (
            .O(N__36608),
            .I(N__36605));
    LocalMux I__7611 (
            .O(N__36605),
            .I(N__36602));
    Span4Mux_s2_v I__7610 (
            .O(N__36602),
            .I(N__36599));
    Span4Mux_v I__7609 (
            .O(N__36599),
            .I(N__36595));
    InMux I__7608 (
            .O(N__36598),
            .I(N__36592));
    Odrv4 I__7607 (
            .O(N__36595),
            .I(T01_c));
    LocalMux I__7606 (
            .O(N__36592),
            .I(T01_c));
    InMux I__7605 (
            .O(N__36587),
            .I(N__36583));
    InMux I__7604 (
            .O(N__36586),
            .I(N__36580));
    LocalMux I__7603 (
            .O(N__36583),
            .I(N__36571));
    LocalMux I__7602 (
            .O(N__36580),
            .I(N__36571));
    InMux I__7601 (
            .O(N__36579),
            .I(N__36568));
    InMux I__7600 (
            .O(N__36578),
            .I(N__36565));
    InMux I__7599 (
            .O(N__36577),
            .I(N__36560));
    InMux I__7598 (
            .O(N__36576),
            .I(N__36560));
    Span4Mux_v I__7597 (
            .O(N__36571),
            .I(N__36555));
    LocalMux I__7596 (
            .O(N__36568),
            .I(N__36555));
    LocalMux I__7595 (
            .O(N__36565),
            .I(N__36552));
    LocalMux I__7594 (
            .O(N__36560),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__7593 (
            .O(N__36555),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv4 I__7592 (
            .O(N__36552),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__7591 (
            .O(N__36545),
            .I(N__36542));
    LocalMux I__7590 (
            .O(N__36542),
            .I(N__36539));
    Span4Mux_s2_v I__7589 (
            .O(N__36539),
            .I(N__36536));
    Span4Mux_v I__7588 (
            .O(N__36536),
            .I(N__36532));
    InMux I__7587 (
            .O(N__36535),
            .I(N__36529));
    Odrv4 I__7586 (
            .O(N__36532),
            .I(T23_c));
    LocalMux I__7585 (
            .O(N__36529),
            .I(T23_c));
    InMux I__7584 (
            .O(N__36524),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__7583 (
            .O(N__36521),
            .I(bfn_15_20_0_));
    InMux I__7582 (
            .O(N__36518),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__7581 (
            .O(N__36515),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__7580 (
            .O(N__36512),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    InMux I__7579 (
            .O(N__36509),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__7578 (
            .O(N__36506),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__7577 (
            .O(N__36503),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    InMux I__7576 (
            .O(N__36500),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    InMux I__7575 (
            .O(N__36497),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__7574 (
            .O(N__36494),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    InMux I__7573 (
            .O(N__36491),
            .I(bfn_15_19_0_));
    InMux I__7572 (
            .O(N__36488),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    InMux I__7571 (
            .O(N__36485),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__7570 (
            .O(N__36482),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__7569 (
            .O(N__36479),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__7568 (
            .O(N__36476),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    InMux I__7567 (
            .O(N__36473),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__7566 (
            .O(N__36470),
            .I(N__36467));
    LocalMux I__7565 (
            .O(N__36467),
            .I(N__36464));
    Span4Mux_v I__7564 (
            .O(N__36464),
            .I(N__36461));
    Odrv4 I__7563 (
            .O(N__36461),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__7562 (
            .O(N__36458),
            .I(N__36455));
    LocalMux I__7561 (
            .O(N__36455),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__7560 (
            .O(N__36452),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__7559 (
            .O(N__36449),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__7558 (
            .O(N__36446),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__7557 (
            .O(N__36443),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__7556 (
            .O(N__36440),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__7555 (
            .O(N__36437),
            .I(N__36434));
    InMux I__7554 (
            .O(N__36434),
            .I(N__36431));
    LocalMux I__7553 (
            .O(N__36431),
            .I(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ));
    InMux I__7552 (
            .O(N__36428),
            .I(N__36425));
    LocalMux I__7551 (
            .O(N__36425),
            .I(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ));
    CascadeMux I__7550 (
            .O(N__36422),
            .I(N__36419));
    InMux I__7549 (
            .O(N__36419),
            .I(N__36416));
    LocalMux I__7548 (
            .O(N__36416),
            .I(N__36413));
    Odrv4 I__7547 (
            .O(N__36413),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    CascadeMux I__7546 (
            .O(N__36410),
            .I(N__36407));
    InMux I__7545 (
            .O(N__36407),
            .I(N__36404));
    LocalMux I__7544 (
            .O(N__36404),
            .I(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ));
    CascadeMux I__7543 (
            .O(N__36401),
            .I(N__36398));
    InMux I__7542 (
            .O(N__36398),
            .I(N__36395));
    LocalMux I__7541 (
            .O(N__36395),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__7540 (
            .O(N__36392),
            .I(N__36389));
    LocalMux I__7539 (
            .O(N__36389),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    CascadeMux I__7538 (
            .O(N__36386),
            .I(N__36383));
    InMux I__7537 (
            .O(N__36383),
            .I(N__36380));
    LocalMux I__7536 (
            .O(N__36380),
            .I(N__36377));
    Odrv4 I__7535 (
            .O(N__36377),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    CascadeMux I__7534 (
            .O(N__36374),
            .I(N__36371));
    InMux I__7533 (
            .O(N__36371),
            .I(N__36368));
    LocalMux I__7532 (
            .O(N__36368),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__7531 (
            .O(N__36365),
            .I(N__36362));
    LocalMux I__7530 (
            .O(N__36362),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    CascadeMux I__7529 (
            .O(N__36359),
            .I(N__36356));
    InMux I__7528 (
            .O(N__36356),
            .I(N__36353));
    LocalMux I__7527 (
            .O(N__36353),
            .I(N__36350));
    Span4Mux_h I__7526 (
            .O(N__36350),
            .I(N__36347));
    Odrv4 I__7525 (
            .O(N__36347),
            .I(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ));
    InMux I__7524 (
            .O(N__36344),
            .I(N__36341));
    LocalMux I__7523 (
            .O(N__36341),
            .I(N__36338));
    Odrv4 I__7522 (
            .O(N__36338),
            .I(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ));
    CascadeMux I__7521 (
            .O(N__36335),
            .I(N__36332));
    InMux I__7520 (
            .O(N__36332),
            .I(N__36329));
    LocalMux I__7519 (
            .O(N__36329),
            .I(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ));
    InMux I__7518 (
            .O(N__36326),
            .I(N__36323));
    LocalMux I__7517 (
            .O(N__36323),
            .I(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ));
    InMux I__7516 (
            .O(N__36320),
            .I(N__36317));
    LocalMux I__7515 (
            .O(N__36317),
            .I(N__36314));
    Odrv4 I__7514 (
            .O(N__36314),
            .I(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ));
    CascadeMux I__7513 (
            .O(N__36311),
            .I(N__36308));
    InMux I__7512 (
            .O(N__36308),
            .I(N__36305));
    LocalMux I__7511 (
            .O(N__36305),
            .I(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ));
    InMux I__7510 (
            .O(N__36302),
            .I(N__36299));
    LocalMux I__7509 (
            .O(N__36299),
            .I(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ));
    CascadeMux I__7508 (
            .O(N__36296),
            .I(N__36293));
    InMux I__7507 (
            .O(N__36293),
            .I(N__36290));
    LocalMux I__7506 (
            .O(N__36290),
            .I(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ));
    CascadeMux I__7505 (
            .O(N__36287),
            .I(N__36283));
    InMux I__7504 (
            .O(N__36286),
            .I(N__36280));
    InMux I__7503 (
            .O(N__36283),
            .I(N__36276));
    LocalMux I__7502 (
            .O(N__36280),
            .I(N__36273));
    InMux I__7501 (
            .O(N__36279),
            .I(N__36270));
    LocalMux I__7500 (
            .O(N__36276),
            .I(N__36267));
    Span4Mux_v I__7499 (
            .O(N__36273),
            .I(N__36264));
    LocalMux I__7498 (
            .O(N__36270),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__7497 (
            .O(N__36267),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    Odrv4 I__7496 (
            .O(N__36264),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__7495 (
            .O(N__36257),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__7494 (
            .O(N__36254),
            .I(N__36250));
    InMux I__7493 (
            .O(N__36253),
            .I(N__36247));
    LocalMux I__7492 (
            .O(N__36250),
            .I(N__36244));
    LocalMux I__7491 (
            .O(N__36247),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    Odrv12 I__7490 (
            .O(N__36244),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__7489 (
            .O(N__36239),
            .I(N__36236));
    InMux I__7488 (
            .O(N__36236),
            .I(N__36231));
    InMux I__7487 (
            .O(N__36235),
            .I(N__36228));
    InMux I__7486 (
            .O(N__36234),
            .I(N__36225));
    LocalMux I__7485 (
            .O(N__36231),
            .I(N__36218));
    LocalMux I__7484 (
            .O(N__36228),
            .I(N__36218));
    LocalMux I__7483 (
            .O(N__36225),
            .I(N__36218));
    Odrv4 I__7482 (
            .O(N__36218),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__7481 (
            .O(N__36215),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__7480 (
            .O(N__36212),
            .I(N__36208));
    InMux I__7479 (
            .O(N__36211),
            .I(N__36205));
    LocalMux I__7478 (
            .O(N__36208),
            .I(N__36202));
    LocalMux I__7477 (
            .O(N__36205),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    Odrv12 I__7476 (
            .O(N__36202),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__7475 (
            .O(N__36197),
            .I(N__36194));
    InMux I__7474 (
            .O(N__36194),
            .I(N__36189));
    InMux I__7473 (
            .O(N__36193),
            .I(N__36186));
    InMux I__7472 (
            .O(N__36192),
            .I(N__36183));
    LocalMux I__7471 (
            .O(N__36189),
            .I(N__36178));
    LocalMux I__7470 (
            .O(N__36186),
            .I(N__36178));
    LocalMux I__7469 (
            .O(N__36183),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    Odrv4 I__7468 (
            .O(N__36178),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__7467 (
            .O(N__36173),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__7466 (
            .O(N__36170),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__7465 (
            .O(N__36167),
            .I(N__36163));
    CEMux I__7464 (
            .O(N__36166),
            .I(N__36160));
    LocalMux I__7463 (
            .O(N__36163),
            .I(N__36154));
    LocalMux I__7462 (
            .O(N__36160),
            .I(N__36151));
    CEMux I__7461 (
            .O(N__36159),
            .I(N__36148));
    CEMux I__7460 (
            .O(N__36158),
            .I(N__36145));
    CEMux I__7459 (
            .O(N__36157),
            .I(N__36142));
    Span4Mux_v I__7458 (
            .O(N__36154),
            .I(N__36139));
    Span4Mux_v I__7457 (
            .O(N__36151),
            .I(N__36136));
    LocalMux I__7456 (
            .O(N__36148),
            .I(N__36133));
    LocalMux I__7455 (
            .O(N__36145),
            .I(N__36130));
    LocalMux I__7454 (
            .O(N__36142),
            .I(N__36127));
    Span4Mux_h I__7453 (
            .O(N__36139),
            .I(N__36124));
    Span4Mux_h I__7452 (
            .O(N__36136),
            .I(N__36119));
    Span4Mux_h I__7451 (
            .O(N__36133),
            .I(N__36119));
    Span4Mux_v I__7450 (
            .O(N__36130),
            .I(N__36116));
    Span4Mux_h I__7449 (
            .O(N__36127),
            .I(N__36113));
    Span4Mux_v I__7448 (
            .O(N__36124),
            .I(N__36108));
    Span4Mux_h I__7447 (
            .O(N__36119),
            .I(N__36108));
    Span4Mux_h I__7446 (
            .O(N__36116),
            .I(N__36103));
    Span4Mux_h I__7445 (
            .O(N__36113),
            .I(N__36103));
    Odrv4 I__7444 (
            .O(N__36108),
            .I(\delay_measurement_inst.delay_tr_timer.N_204_i ));
    Odrv4 I__7443 (
            .O(N__36103),
            .I(\delay_measurement_inst.delay_tr_timer.N_204_i ));
    InMux I__7442 (
            .O(N__36098),
            .I(N__36095));
    LocalMux I__7441 (
            .O(N__36095),
            .I(N__36092));
    Span4Mux_h I__7440 (
            .O(N__36092),
            .I(N__36089));
    Odrv4 I__7439 (
            .O(N__36089),
            .I(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ));
    CascadeMux I__7438 (
            .O(N__36086),
            .I(N__36083));
    InMux I__7437 (
            .O(N__36083),
            .I(N__36080));
    LocalMux I__7436 (
            .O(N__36080),
            .I(N__36077));
    Odrv4 I__7435 (
            .O(N__36077),
            .I(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ));
    InMux I__7434 (
            .O(N__36074),
            .I(N__36071));
    LocalMux I__7433 (
            .O(N__36071),
            .I(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ));
    CascadeMux I__7432 (
            .O(N__36068),
            .I(N__36065));
    InMux I__7431 (
            .O(N__36065),
            .I(N__36062));
    LocalMux I__7430 (
            .O(N__36062),
            .I(N__36059));
    Span4Mux_v I__7429 (
            .O(N__36059),
            .I(N__36056));
    Odrv4 I__7428 (
            .O(N__36056),
            .I(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ));
    InMux I__7427 (
            .O(N__36053),
            .I(N__36050));
    LocalMux I__7426 (
            .O(N__36050),
            .I(N__36047));
    Sp12to4 I__7425 (
            .O(N__36047),
            .I(N__36044));
    Odrv12 I__7424 (
            .O(N__36044),
            .I(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ));
    CascadeMux I__7423 (
            .O(N__36041),
            .I(N__36037));
    CascadeMux I__7422 (
            .O(N__36040),
            .I(N__36034));
    InMux I__7421 (
            .O(N__36037),
            .I(N__36031));
    InMux I__7420 (
            .O(N__36034),
            .I(N__36027));
    LocalMux I__7419 (
            .O(N__36031),
            .I(N__36024));
    InMux I__7418 (
            .O(N__36030),
            .I(N__36021));
    LocalMux I__7417 (
            .O(N__36027),
            .I(N__36018));
    Span4Mux_v I__7416 (
            .O(N__36024),
            .I(N__36015));
    LocalMux I__7415 (
            .O(N__36021),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__7414 (
            .O(N__36018),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    Odrv4 I__7413 (
            .O(N__36015),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__7412 (
            .O(N__36008),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__7411 (
            .O(N__36005),
            .I(N__36002));
    InMux I__7410 (
            .O(N__36002),
            .I(N__35997));
    InMux I__7409 (
            .O(N__36001),
            .I(N__35994));
    InMux I__7408 (
            .O(N__36000),
            .I(N__35991));
    LocalMux I__7407 (
            .O(N__35997),
            .I(N__35984));
    LocalMux I__7406 (
            .O(N__35994),
            .I(N__35984));
    LocalMux I__7405 (
            .O(N__35991),
            .I(N__35984));
    Odrv4 I__7404 (
            .O(N__35984),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__7403 (
            .O(N__35981),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__7402 (
            .O(N__35978),
            .I(N__35971));
    InMux I__7401 (
            .O(N__35977),
            .I(N__35971));
    InMux I__7400 (
            .O(N__35976),
            .I(N__35968));
    LocalMux I__7399 (
            .O(N__35971),
            .I(N__35965));
    LocalMux I__7398 (
            .O(N__35968),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    Odrv4 I__7397 (
            .O(N__35965),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__7396 (
            .O(N__35960),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__7395 (
            .O(N__35957),
            .I(N__35950));
    InMux I__7394 (
            .O(N__35956),
            .I(N__35950));
    InMux I__7393 (
            .O(N__35955),
            .I(N__35947));
    LocalMux I__7392 (
            .O(N__35950),
            .I(N__35944));
    LocalMux I__7391 (
            .O(N__35947),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    Odrv4 I__7390 (
            .O(N__35944),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__7389 (
            .O(N__35939),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__7388 (
            .O(N__35936),
            .I(N__35932));
    InMux I__7387 (
            .O(N__35935),
            .I(N__35928));
    InMux I__7386 (
            .O(N__35932),
            .I(N__35925));
    InMux I__7385 (
            .O(N__35931),
            .I(N__35922));
    LocalMux I__7384 (
            .O(N__35928),
            .I(N__35917));
    LocalMux I__7383 (
            .O(N__35925),
            .I(N__35917));
    LocalMux I__7382 (
            .O(N__35922),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    Odrv12 I__7381 (
            .O(N__35917),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__7380 (
            .O(N__35912),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__7379 (
            .O(N__35909),
            .I(N__35905));
    CascadeMux I__7378 (
            .O(N__35908),
            .I(N__35902));
    InMux I__7377 (
            .O(N__35905),
            .I(N__35896));
    InMux I__7376 (
            .O(N__35902),
            .I(N__35896));
    InMux I__7375 (
            .O(N__35901),
            .I(N__35893));
    LocalMux I__7374 (
            .O(N__35896),
            .I(N__35890));
    LocalMux I__7373 (
            .O(N__35893),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    Odrv12 I__7372 (
            .O(N__35890),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__7371 (
            .O(N__35885),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__7370 (
            .O(N__35882),
            .I(N__35878));
    CascadeMux I__7369 (
            .O(N__35881),
            .I(N__35875));
    InMux I__7368 (
            .O(N__35878),
            .I(N__35869));
    InMux I__7367 (
            .O(N__35875),
            .I(N__35869));
    InMux I__7366 (
            .O(N__35874),
            .I(N__35866));
    LocalMux I__7365 (
            .O(N__35869),
            .I(N__35863));
    LocalMux I__7364 (
            .O(N__35866),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    Odrv4 I__7363 (
            .O(N__35863),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__7362 (
            .O(N__35858),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__7361 (
            .O(N__35855),
            .I(N__35852));
    InMux I__7360 (
            .O(N__35852),
            .I(N__35848));
    InMux I__7359 (
            .O(N__35851),
            .I(N__35845));
    LocalMux I__7358 (
            .O(N__35848),
            .I(N__35839));
    LocalMux I__7357 (
            .O(N__35845),
            .I(N__35839));
    InMux I__7356 (
            .O(N__35844),
            .I(N__35836));
    Span4Mux_v I__7355 (
            .O(N__35839),
            .I(N__35833));
    LocalMux I__7354 (
            .O(N__35836),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    Odrv4 I__7353 (
            .O(N__35833),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__7352 (
            .O(N__35828),
            .I(bfn_15_13_0_));
    CascadeMux I__7351 (
            .O(N__35825),
            .I(N__35820));
    InMux I__7350 (
            .O(N__35824),
            .I(N__35817));
    InMux I__7349 (
            .O(N__35823),
            .I(N__35814));
    InMux I__7348 (
            .O(N__35820),
            .I(N__35811));
    LocalMux I__7347 (
            .O(N__35817),
            .I(N__35808));
    LocalMux I__7346 (
            .O(N__35814),
            .I(N__35801));
    LocalMux I__7345 (
            .O(N__35811),
            .I(N__35801));
    Span4Mux_v I__7344 (
            .O(N__35808),
            .I(N__35801));
    Odrv4 I__7343 (
            .O(N__35801),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__7342 (
            .O(N__35798),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__7341 (
            .O(N__35795),
            .I(N__35788));
    InMux I__7340 (
            .O(N__35794),
            .I(N__35788));
    InMux I__7339 (
            .O(N__35793),
            .I(N__35785));
    LocalMux I__7338 (
            .O(N__35788),
            .I(N__35782));
    LocalMux I__7337 (
            .O(N__35785),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    Odrv4 I__7336 (
            .O(N__35782),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__7335 (
            .O(N__35777),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__7334 (
            .O(N__35774),
            .I(N__35771));
    InMux I__7333 (
            .O(N__35771),
            .I(N__35766));
    InMux I__7332 (
            .O(N__35770),
            .I(N__35763));
    InMux I__7331 (
            .O(N__35769),
            .I(N__35760));
    LocalMux I__7330 (
            .O(N__35766),
            .I(N__35755));
    LocalMux I__7329 (
            .O(N__35763),
            .I(N__35755));
    LocalMux I__7328 (
            .O(N__35760),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    Odrv12 I__7327 (
            .O(N__35755),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__7326 (
            .O(N__35750),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__7325 (
            .O(N__35747),
            .I(N__35743));
    CascadeMux I__7324 (
            .O(N__35746),
            .I(N__35740));
    InMux I__7323 (
            .O(N__35743),
            .I(N__35734));
    InMux I__7322 (
            .O(N__35740),
            .I(N__35734));
    InMux I__7321 (
            .O(N__35739),
            .I(N__35731));
    LocalMux I__7320 (
            .O(N__35734),
            .I(N__35728));
    LocalMux I__7319 (
            .O(N__35731),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    Odrv12 I__7318 (
            .O(N__35728),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__7317 (
            .O(N__35723),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__7316 (
            .O(N__35720),
            .I(N__35717));
    InMux I__7315 (
            .O(N__35717),
            .I(N__35712));
    InMux I__7314 (
            .O(N__35716),
            .I(N__35709));
    InMux I__7313 (
            .O(N__35715),
            .I(N__35706));
    LocalMux I__7312 (
            .O(N__35712),
            .I(N__35701));
    LocalMux I__7311 (
            .O(N__35709),
            .I(N__35701));
    LocalMux I__7310 (
            .O(N__35706),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    Odrv12 I__7309 (
            .O(N__35701),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__7308 (
            .O(N__35696),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__7307 (
            .O(N__35693),
            .I(N__35690));
    InMux I__7306 (
            .O(N__35690),
            .I(N__35685));
    InMux I__7305 (
            .O(N__35689),
            .I(N__35682));
    InMux I__7304 (
            .O(N__35688),
            .I(N__35679));
    LocalMux I__7303 (
            .O(N__35685),
            .I(N__35674));
    LocalMux I__7302 (
            .O(N__35682),
            .I(N__35674));
    LocalMux I__7301 (
            .O(N__35679),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    Odrv12 I__7300 (
            .O(N__35674),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__7299 (
            .O(N__35669),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__7298 (
            .O(N__35666),
            .I(N__35661));
    InMux I__7297 (
            .O(N__35665),
            .I(N__35656));
    InMux I__7296 (
            .O(N__35664),
            .I(N__35656));
    LocalMux I__7295 (
            .O(N__35661),
            .I(N__35651));
    LocalMux I__7294 (
            .O(N__35656),
            .I(N__35651));
    Odrv4 I__7293 (
            .O(N__35651),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__7292 (
            .O(N__35648),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__7291 (
            .O(N__35645),
            .I(N__35641));
    InMux I__7290 (
            .O(N__35644),
            .I(N__35638));
    InMux I__7289 (
            .O(N__35641),
            .I(N__35634));
    LocalMux I__7288 (
            .O(N__35638),
            .I(N__35631));
    InMux I__7287 (
            .O(N__35637),
            .I(N__35628));
    LocalMux I__7286 (
            .O(N__35634),
            .I(N__35623));
    Span4Mux_v I__7285 (
            .O(N__35631),
            .I(N__35623));
    LocalMux I__7284 (
            .O(N__35628),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    Odrv4 I__7283 (
            .O(N__35623),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__7282 (
            .O(N__35618),
            .I(bfn_15_12_0_));
    InMux I__7281 (
            .O(N__35615),
            .I(N__35612));
    LocalMux I__7280 (
            .O(N__35612),
            .I(N__35608));
    InMux I__7279 (
            .O(N__35611),
            .I(N__35605));
    Span4Mux_h I__7278 (
            .O(N__35608),
            .I(N__35601));
    LocalMux I__7277 (
            .O(N__35605),
            .I(N__35598));
    InMux I__7276 (
            .O(N__35604),
            .I(N__35595));
    Odrv4 I__7275 (
            .O(N__35601),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    Odrv4 I__7274 (
            .O(N__35598),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__7273 (
            .O(N__35595),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__7272 (
            .O(N__35588),
            .I(N__35584));
    CascadeMux I__7271 (
            .O(N__35587),
            .I(N__35581));
    LocalMux I__7270 (
            .O(N__35584),
            .I(N__35578));
    InMux I__7269 (
            .O(N__35581),
            .I(N__35574));
    Span4Mux_h I__7268 (
            .O(N__35578),
            .I(N__35571));
    InMux I__7267 (
            .O(N__35577),
            .I(N__35568));
    LocalMux I__7266 (
            .O(N__35574),
            .I(N__35565));
    Odrv4 I__7265 (
            .O(N__35571),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__7264 (
            .O(N__35568),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    Odrv12 I__7263 (
            .O(N__35565),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__7262 (
            .O(N__35558),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__7261 (
            .O(N__35555),
            .I(N__35551));
    CascadeMux I__7260 (
            .O(N__35554),
            .I(N__35548));
    InMux I__7259 (
            .O(N__35551),
            .I(N__35542));
    InMux I__7258 (
            .O(N__35548),
            .I(N__35542));
    InMux I__7257 (
            .O(N__35547),
            .I(N__35539));
    LocalMux I__7256 (
            .O(N__35542),
            .I(N__35536));
    LocalMux I__7255 (
            .O(N__35539),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    Odrv12 I__7254 (
            .O(N__35536),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__7253 (
            .O(N__35531),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__7252 (
            .O(N__35528),
            .I(N__35521));
    InMux I__7251 (
            .O(N__35527),
            .I(N__35521));
    InMux I__7250 (
            .O(N__35526),
            .I(N__35518));
    LocalMux I__7249 (
            .O(N__35521),
            .I(N__35515));
    LocalMux I__7248 (
            .O(N__35518),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    Odrv4 I__7247 (
            .O(N__35515),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__7246 (
            .O(N__35510),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__7245 (
            .O(N__35507),
            .I(N__35504));
    InMux I__7244 (
            .O(N__35504),
            .I(N__35499));
    InMux I__7243 (
            .O(N__35503),
            .I(N__35496));
    InMux I__7242 (
            .O(N__35502),
            .I(N__35493));
    LocalMux I__7241 (
            .O(N__35499),
            .I(N__35488));
    LocalMux I__7240 (
            .O(N__35496),
            .I(N__35488));
    LocalMux I__7239 (
            .O(N__35493),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    Odrv12 I__7238 (
            .O(N__35488),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__7237 (
            .O(N__35483),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__7236 (
            .O(N__35480),
            .I(N__35476));
    CascadeMux I__7235 (
            .O(N__35479),
            .I(N__35473));
    InMux I__7234 (
            .O(N__35476),
            .I(N__35467));
    InMux I__7233 (
            .O(N__35473),
            .I(N__35467));
    InMux I__7232 (
            .O(N__35472),
            .I(N__35464));
    LocalMux I__7231 (
            .O(N__35467),
            .I(N__35461));
    LocalMux I__7230 (
            .O(N__35464),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    Odrv4 I__7229 (
            .O(N__35461),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__7228 (
            .O(N__35456),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__7227 (
            .O(N__35453),
            .I(N__35448));
    InMux I__7226 (
            .O(N__35452),
            .I(N__35443));
    InMux I__7225 (
            .O(N__35451),
            .I(N__35443));
    LocalMux I__7224 (
            .O(N__35448),
            .I(N__35438));
    LocalMux I__7223 (
            .O(N__35443),
            .I(N__35438));
    Odrv4 I__7222 (
            .O(N__35438),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__7221 (
            .O(N__35435),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__7220 (
            .O(N__35432),
            .I(N__35429));
    InMux I__7219 (
            .O(N__35429),
            .I(N__35424));
    InMux I__7218 (
            .O(N__35428),
            .I(N__35421));
    InMux I__7217 (
            .O(N__35427),
            .I(N__35418));
    LocalMux I__7216 (
            .O(N__35424),
            .I(N__35413));
    LocalMux I__7215 (
            .O(N__35421),
            .I(N__35413));
    LocalMux I__7214 (
            .O(N__35418),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    Odrv12 I__7213 (
            .O(N__35413),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__7212 (
            .O(N__35408),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__7211 (
            .O(N__35405),
            .I(N__35401));
    CascadeMux I__7210 (
            .O(N__35404),
            .I(N__35398));
    InMux I__7209 (
            .O(N__35401),
            .I(N__35395));
    InMux I__7208 (
            .O(N__35398),
            .I(N__35391));
    LocalMux I__7207 (
            .O(N__35395),
            .I(N__35388));
    InMux I__7206 (
            .O(N__35394),
            .I(N__35385));
    LocalMux I__7205 (
            .O(N__35391),
            .I(N__35382));
    Span4Mux_v I__7204 (
            .O(N__35388),
            .I(N__35379));
    LocalMux I__7203 (
            .O(N__35385),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__7202 (
            .O(N__35382),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    Odrv4 I__7201 (
            .O(N__35379),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__7200 (
            .O(N__35372),
            .I(bfn_15_11_0_));
    InMux I__7199 (
            .O(N__35369),
            .I(N__35366));
    LocalMux I__7198 (
            .O(N__35366),
            .I(N__35363));
    Odrv4 I__7197 (
            .O(N__35363),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    CascadeMux I__7196 (
            .O(N__35360),
            .I(N__35357));
    InMux I__7195 (
            .O(N__35357),
            .I(N__35354));
    LocalMux I__7194 (
            .O(N__35354),
            .I(N__35351));
    Span4Mux_v I__7193 (
            .O(N__35351),
            .I(N__35348));
    Odrv4 I__7192 (
            .O(N__35348),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    InMux I__7191 (
            .O(N__35345),
            .I(N__35342));
    LocalMux I__7190 (
            .O(N__35342),
            .I(N__35339));
    Odrv4 I__7189 (
            .O(N__35339),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    CascadeMux I__7188 (
            .O(N__35336),
            .I(N__35333));
    InMux I__7187 (
            .O(N__35333),
            .I(N__35329));
    InMux I__7186 (
            .O(N__35332),
            .I(N__35326));
    LocalMux I__7185 (
            .O(N__35329),
            .I(N__35323));
    LocalMux I__7184 (
            .O(N__35326),
            .I(N__35320));
    Odrv4 I__7183 (
            .O(N__35323),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    Odrv4 I__7182 (
            .O(N__35320),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    InMux I__7181 (
            .O(N__35315),
            .I(N__35312));
    LocalMux I__7180 (
            .O(N__35312),
            .I(N__35309));
    Span4Mux_h I__7179 (
            .O(N__35309),
            .I(N__35306));
    Odrv4 I__7178 (
            .O(N__35306),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ));
    InMux I__7177 (
            .O(N__35303),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ));
    InMux I__7176 (
            .O(N__35300),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ));
    InMux I__7175 (
            .O(N__35297),
            .I(N__35293));
    InMux I__7174 (
            .O(N__35296),
            .I(N__35290));
    LocalMux I__7173 (
            .O(N__35293),
            .I(N__35287));
    LocalMux I__7172 (
            .O(N__35290),
            .I(N__35284));
    Span4Mux_h I__7171 (
            .O(N__35287),
            .I(N__35281));
    Span4Mux_h I__7170 (
            .O(N__35284),
            .I(N__35278));
    Odrv4 I__7169 (
            .O(N__35281),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    Odrv4 I__7168 (
            .O(N__35278),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ));
    InMux I__7167 (
            .O(N__35273),
            .I(N__35269));
    InMux I__7166 (
            .O(N__35272),
            .I(N__35266));
    LocalMux I__7165 (
            .O(N__35269),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    LocalMux I__7164 (
            .O(N__35266),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__7163 (
            .O(N__35261),
            .I(N__35258));
    LocalMux I__7162 (
            .O(N__35258),
            .I(N__35255));
    Odrv4 I__7161 (
            .O(N__35255),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__7160 (
            .O(N__35252),
            .I(N__35248));
    InMux I__7159 (
            .O(N__35251),
            .I(N__35245));
    LocalMux I__7158 (
            .O(N__35248),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    LocalMux I__7157 (
            .O(N__35245),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    CascadeMux I__7156 (
            .O(N__35240),
            .I(N__35237));
    InMux I__7155 (
            .O(N__35237),
            .I(N__35234));
    LocalMux I__7154 (
            .O(N__35234),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__7153 (
            .O(N__35231),
            .I(N__35227));
    InMux I__7152 (
            .O(N__35230),
            .I(N__35224));
    LocalMux I__7151 (
            .O(N__35227),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    LocalMux I__7150 (
            .O(N__35224),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__7149 (
            .O(N__35219),
            .I(N__35216));
    LocalMux I__7148 (
            .O(N__35216),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__7147 (
            .O(N__35213),
            .I(N__35209));
    InMux I__7146 (
            .O(N__35212),
            .I(N__35206));
    LocalMux I__7145 (
            .O(N__35209),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    LocalMux I__7144 (
            .O(N__35206),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__7143 (
            .O(N__35201),
            .I(N__35198));
    LocalMux I__7142 (
            .O(N__35198),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__7141 (
            .O(N__35195),
            .I(N__35192));
    LocalMux I__7140 (
            .O(N__35192),
            .I(N__35189));
    Span4Mux_h I__7139 (
            .O(N__35189),
            .I(N__35186));
    Odrv4 I__7138 (
            .O(N__35186),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    InMux I__7137 (
            .O(N__35183),
            .I(N__35179));
    InMux I__7136 (
            .O(N__35182),
            .I(N__35176));
    LocalMux I__7135 (
            .O(N__35179),
            .I(N__35173));
    LocalMux I__7134 (
            .O(N__35176),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__7133 (
            .O(N__35173),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    CascadeMux I__7132 (
            .O(N__35168),
            .I(N__35165));
    InMux I__7131 (
            .O(N__35165),
            .I(N__35162));
    LocalMux I__7130 (
            .O(N__35162),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    InMux I__7129 (
            .O(N__35159),
            .I(N__35156));
    LocalMux I__7128 (
            .O(N__35156),
            .I(N__35153));
    Span4Mux_h I__7127 (
            .O(N__35153),
            .I(N__35150));
    Span4Mux_h I__7126 (
            .O(N__35150),
            .I(N__35147));
    Odrv4 I__7125 (
            .O(N__35147),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    InMux I__7124 (
            .O(N__35144),
            .I(N__35140));
    InMux I__7123 (
            .O(N__35143),
            .I(N__35137));
    LocalMux I__7122 (
            .O(N__35140),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    LocalMux I__7121 (
            .O(N__35137),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    CascadeMux I__7120 (
            .O(N__35132),
            .I(N__35129));
    InMux I__7119 (
            .O(N__35129),
            .I(N__35126));
    LocalMux I__7118 (
            .O(N__35126),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__7117 (
            .O(N__35123),
            .I(N__35120));
    LocalMux I__7116 (
            .O(N__35120),
            .I(N__35117));
    Odrv4 I__7115 (
            .O(N__35117),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    InMux I__7114 (
            .O(N__35114),
            .I(N__35110));
    InMux I__7113 (
            .O(N__35113),
            .I(N__35107));
    LocalMux I__7112 (
            .O(N__35110),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    LocalMux I__7111 (
            .O(N__35107),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    CascadeMux I__7110 (
            .O(N__35102),
            .I(N__35099));
    InMux I__7109 (
            .O(N__35099),
            .I(N__35096));
    LocalMux I__7108 (
            .O(N__35096),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__7107 (
            .O(N__35093),
            .I(N__35090));
    LocalMux I__7106 (
            .O(N__35090),
            .I(N__35087));
    Odrv4 I__7105 (
            .O(N__35087),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    CascadeMux I__7104 (
            .O(N__35084),
            .I(N__35081));
    InMux I__7103 (
            .O(N__35081),
            .I(N__35078));
    LocalMux I__7102 (
            .O(N__35078),
            .I(N__35075));
    Odrv12 I__7101 (
            .O(N__35075),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    InMux I__7100 (
            .O(N__35072),
            .I(N__35068));
    InMux I__7099 (
            .O(N__35071),
            .I(N__35065));
    LocalMux I__7098 (
            .O(N__35068),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    LocalMux I__7097 (
            .O(N__35065),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__7096 (
            .O(N__35060),
            .I(N__35057));
    LocalMux I__7095 (
            .O(N__35057),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__7094 (
            .O(N__35054),
            .I(N__35051));
    InMux I__7093 (
            .O(N__35051),
            .I(N__35048));
    LocalMux I__7092 (
            .O(N__35048),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__7091 (
            .O(N__35045),
            .I(N__35041));
    InMux I__7090 (
            .O(N__35044),
            .I(N__35038));
    LocalMux I__7089 (
            .O(N__35041),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    LocalMux I__7088 (
            .O(N__35038),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    CascadeMux I__7087 (
            .O(N__35033),
            .I(N__35030));
    InMux I__7086 (
            .O(N__35030),
            .I(N__35027));
    LocalMux I__7085 (
            .O(N__35027),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__7084 (
            .O(N__35024),
            .I(N__35021));
    LocalMux I__7083 (
            .O(N__35021),
            .I(N__35018));
    Odrv4 I__7082 (
            .O(N__35018),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    InMux I__7081 (
            .O(N__35015),
            .I(N__35011));
    InMux I__7080 (
            .O(N__35014),
            .I(N__35008));
    LocalMux I__7079 (
            .O(N__35011),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    LocalMux I__7078 (
            .O(N__35008),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    CascadeMux I__7077 (
            .O(N__35003),
            .I(N__35000));
    InMux I__7076 (
            .O(N__35000),
            .I(N__34997));
    LocalMux I__7075 (
            .O(N__34997),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__7074 (
            .O(N__34994),
            .I(N__34991));
    LocalMux I__7073 (
            .O(N__34991),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    InMux I__7072 (
            .O(N__34988),
            .I(N__34984));
    InMux I__7071 (
            .O(N__34987),
            .I(N__34981));
    LocalMux I__7070 (
            .O(N__34984),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    LocalMux I__7069 (
            .O(N__34981),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    CascadeMux I__7068 (
            .O(N__34976),
            .I(N__34973));
    InMux I__7067 (
            .O(N__34973),
            .I(N__34970));
    LocalMux I__7066 (
            .O(N__34970),
            .I(N__34967));
    Odrv4 I__7065 (
            .O(N__34967),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    InMux I__7064 (
            .O(N__34964),
            .I(N__34960));
    InMux I__7063 (
            .O(N__34963),
            .I(N__34957));
    LocalMux I__7062 (
            .O(N__34960),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    LocalMux I__7061 (
            .O(N__34957),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    CascadeMux I__7060 (
            .O(N__34952),
            .I(N__34949));
    InMux I__7059 (
            .O(N__34949),
            .I(N__34946));
    LocalMux I__7058 (
            .O(N__34946),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__7057 (
            .O(N__34943),
            .I(N__34940));
    LocalMux I__7056 (
            .O(N__34940),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    InMux I__7055 (
            .O(N__34937),
            .I(N__34933));
    InMux I__7054 (
            .O(N__34936),
            .I(N__34930));
    LocalMux I__7053 (
            .O(N__34933),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    LocalMux I__7052 (
            .O(N__34930),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    CascadeMux I__7051 (
            .O(N__34925),
            .I(N__34922));
    InMux I__7050 (
            .O(N__34922),
            .I(N__34919));
    LocalMux I__7049 (
            .O(N__34919),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    InMux I__7048 (
            .O(N__34916),
            .I(N__34912));
    InMux I__7047 (
            .O(N__34915),
            .I(N__34909));
    LocalMux I__7046 (
            .O(N__34912),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    LocalMux I__7045 (
            .O(N__34909),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    CascadeMux I__7044 (
            .O(N__34904),
            .I(N__34901));
    InMux I__7043 (
            .O(N__34901),
            .I(N__34898));
    LocalMux I__7042 (
            .O(N__34898),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__7041 (
            .O(N__34895),
            .I(N__34889));
    InMux I__7040 (
            .O(N__34894),
            .I(N__34886));
    InMux I__7039 (
            .O(N__34893),
            .I(N__34883));
    InMux I__7038 (
            .O(N__34892),
            .I(N__34880));
    LocalMux I__7037 (
            .O(N__34889),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__7036 (
            .O(N__34886),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__7035 (
            .O(N__34883),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__7034 (
            .O(N__34880),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    IoInMux I__7033 (
            .O(N__34871),
            .I(N__34868));
    LocalMux I__7032 (
            .O(N__34868),
            .I(N__34865));
    Span4Mux_s1_v I__7031 (
            .O(N__34865),
            .I(N__34862));
    Span4Mux_v I__7030 (
            .O(N__34862),
            .I(N__34857));
    InMux I__7029 (
            .O(N__34861),
            .I(N__34854));
    InMux I__7028 (
            .O(N__34860),
            .I(N__34851));
    Odrv4 I__7027 (
            .O(N__34857),
            .I(s1_phy_c));
    LocalMux I__7026 (
            .O(N__34854),
            .I(s1_phy_c));
    LocalMux I__7025 (
            .O(N__34851),
            .I(s1_phy_c));
    CascadeMux I__7024 (
            .O(N__34844),
            .I(N__34839));
    InMux I__7023 (
            .O(N__34843),
            .I(N__34835));
    InMux I__7022 (
            .O(N__34842),
            .I(N__34832));
    InMux I__7021 (
            .O(N__34839),
            .I(N__34829));
    InMux I__7020 (
            .O(N__34838),
            .I(N__34826));
    LocalMux I__7019 (
            .O(N__34835),
            .I(N__34823));
    LocalMux I__7018 (
            .O(N__34832),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7017 (
            .O(N__34829),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__7016 (
            .O(N__34826),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv4 I__7015 (
            .O(N__34823),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__7014 (
            .O(N__34814),
            .I(N__34811));
    LocalMux I__7013 (
            .O(N__34811),
            .I(N__34808));
    Span12Mux_s3_v I__7012 (
            .O(N__34808),
            .I(N__34805));
    Odrv12 I__7011 (
            .O(N__34805),
            .I(s2_phy_c));
    InMux I__7010 (
            .O(N__34802),
            .I(N__34796));
    InMux I__7009 (
            .O(N__34801),
            .I(N__34796));
    LocalMux I__7008 (
            .O(N__34796),
            .I(N__34792));
    InMux I__7007 (
            .O(N__34795),
            .I(N__34789));
    Span4Mux_h I__7006 (
            .O(N__34792),
            .I(N__34786));
    LocalMux I__7005 (
            .O(N__34789),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__7004 (
            .O(N__34786),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__7003 (
            .O(N__34781),
            .I(N__34777));
    CascadeMux I__7002 (
            .O(N__34780),
            .I(N__34774));
    InMux I__7001 (
            .O(N__34777),
            .I(N__34771));
    InMux I__7000 (
            .O(N__34774),
            .I(N__34768));
    LocalMux I__6999 (
            .O(N__34771),
            .I(N__34762));
    LocalMux I__6998 (
            .O(N__34768),
            .I(N__34762));
    InMux I__6997 (
            .O(N__34767),
            .I(N__34759));
    Span4Mux_h I__6996 (
            .O(N__34762),
            .I(N__34756));
    LocalMux I__6995 (
            .O(N__34759),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv4 I__6994 (
            .O(N__34756),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__6993 (
            .O(N__34751),
            .I(N__34745));
    InMux I__6992 (
            .O(N__34750),
            .I(N__34745));
    LocalMux I__6991 (
            .O(N__34745),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    InMux I__6990 (
            .O(N__34742),
            .I(N__34739));
    LocalMux I__6989 (
            .O(N__34739),
            .I(N__34736));
    Odrv4 I__6988 (
            .O(N__34736),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__6987 (
            .O(N__34733),
            .I(N__34730));
    InMux I__6986 (
            .O(N__34730),
            .I(N__34725));
    InMux I__6985 (
            .O(N__34729),
            .I(N__34722));
    CascadeMux I__6984 (
            .O(N__34728),
            .I(N__34719));
    LocalMux I__6983 (
            .O(N__34725),
            .I(N__34714));
    LocalMux I__6982 (
            .O(N__34722),
            .I(N__34714));
    InMux I__6981 (
            .O(N__34719),
            .I(N__34711));
    Span4Mux_v I__6980 (
            .O(N__34714),
            .I(N__34708));
    LocalMux I__6979 (
            .O(N__34711),
            .I(N__34703));
    Span4Mux_h I__6978 (
            .O(N__34708),
            .I(N__34703));
    Odrv4 I__6977 (
            .O(N__34703),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    CascadeMux I__6976 (
            .O(N__34700),
            .I(N__34697));
    InMux I__6975 (
            .O(N__34697),
            .I(N__34694));
    LocalMux I__6974 (
            .O(N__34694),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    CascadeMux I__6973 (
            .O(N__34691),
            .I(N__34685));
    InMux I__6972 (
            .O(N__34690),
            .I(N__34682));
    InMux I__6971 (
            .O(N__34689),
            .I(N__34677));
    InMux I__6970 (
            .O(N__34688),
            .I(N__34677));
    InMux I__6969 (
            .O(N__34685),
            .I(N__34674));
    LocalMux I__6968 (
            .O(N__34682),
            .I(N__34671));
    LocalMux I__6967 (
            .O(N__34677),
            .I(N__34668));
    LocalMux I__6966 (
            .O(N__34674),
            .I(N__34663));
    Span4Mux_v I__6965 (
            .O(N__34671),
            .I(N__34663));
    Sp12to4 I__6964 (
            .O(N__34668),
            .I(N__34658));
    Span4Mux_v I__6963 (
            .O(N__34663),
            .I(N__34655));
    InMux I__6962 (
            .O(N__34662),
            .I(N__34652));
    InMux I__6961 (
            .O(N__34661),
            .I(N__34649));
    Span12Mux_v I__6960 (
            .O(N__34658),
            .I(N__34642));
    Sp12to4 I__6959 (
            .O(N__34655),
            .I(N__34642));
    LocalMux I__6958 (
            .O(N__34652),
            .I(N__34642));
    LocalMux I__6957 (
            .O(N__34649),
            .I(phase_controller_inst1_state_4));
    Odrv12 I__6956 (
            .O(N__34642),
            .I(phase_controller_inst1_state_4));
    InMux I__6955 (
            .O(N__34637),
            .I(N__34634));
    LocalMux I__6954 (
            .O(N__34634),
            .I(N__34630));
    InMux I__6953 (
            .O(N__34633),
            .I(N__34627));
    Span4Mux_h I__6952 (
            .O(N__34630),
            .I(N__34622));
    LocalMux I__6951 (
            .O(N__34627),
            .I(N__34622));
    Odrv4 I__6950 (
            .O(N__34622),
            .I(\phase_controller_inst1.time_passed_RNIE87F ));
    CascadeMux I__6949 (
            .O(N__34619),
            .I(N__34616));
    InMux I__6948 (
            .O(N__34616),
            .I(N__34611));
    InMux I__6947 (
            .O(N__34615),
            .I(N__34608));
    InMux I__6946 (
            .O(N__34614),
            .I(N__34605));
    LocalMux I__6945 (
            .O(N__34611),
            .I(N__34602));
    LocalMux I__6944 (
            .O(N__34608),
            .I(N__34597));
    LocalMux I__6943 (
            .O(N__34605),
            .I(N__34597));
    Span4Mux_v I__6942 (
            .O(N__34602),
            .I(N__34592));
    Span4Mux_v I__6941 (
            .O(N__34597),
            .I(N__34592));
    Span4Mux_h I__6940 (
            .O(N__34592),
            .I(N__34589));
    Span4Mux_h I__6939 (
            .O(N__34589),
            .I(N__34585));
    InMux I__6938 (
            .O(N__34588),
            .I(N__34582));
    Span4Mux_v I__6937 (
            .O(N__34585),
            .I(N__34579));
    LocalMux I__6936 (
            .O(N__34582),
            .I(\phase_controller_inst1.hc_time_passed ));
    Odrv4 I__6935 (
            .O(N__34579),
            .I(\phase_controller_inst1.hc_time_passed ));
    CascadeMux I__6934 (
            .O(N__34574),
            .I(N__34569));
    CascadeMux I__6933 (
            .O(N__34573),
            .I(N__34566));
    InMux I__6932 (
            .O(N__34572),
            .I(N__34561));
    InMux I__6931 (
            .O(N__34569),
            .I(N__34561));
    InMux I__6930 (
            .O(N__34566),
            .I(N__34558));
    LocalMux I__6929 (
            .O(N__34561),
            .I(N__34555));
    LocalMux I__6928 (
            .O(N__34558),
            .I(N__34552));
    Span4Mux_v I__6927 (
            .O(N__34555),
            .I(N__34547));
    Span4Mux_v I__6926 (
            .O(N__34552),
            .I(N__34547));
    Odrv4 I__6925 (
            .O(N__34547),
            .I(il_min_comp1_D2));
    InMux I__6924 (
            .O(N__34544),
            .I(N__34541));
    LocalMux I__6923 (
            .O(N__34541),
            .I(N__34538));
    Odrv4 I__6922 (
            .O(N__34538),
            .I(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ));
    InMux I__6921 (
            .O(N__34535),
            .I(N__34530));
    InMux I__6920 (
            .O(N__34534),
            .I(N__34526));
    InMux I__6919 (
            .O(N__34533),
            .I(N__34523));
    LocalMux I__6918 (
            .O(N__34530),
            .I(N__34520));
    InMux I__6917 (
            .O(N__34529),
            .I(N__34517));
    LocalMux I__6916 (
            .O(N__34526),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__6915 (
            .O(N__34523),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__6914 (
            .O(N__34520),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    LocalMux I__6913 (
            .O(N__34517),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__6912 (
            .O(N__34508),
            .I(N__34505));
    LocalMux I__6911 (
            .O(N__34505),
            .I(N__34502));
    Odrv4 I__6910 (
            .O(N__34502),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__6909 (
            .O(N__34499),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__6908 (
            .O(N__34496),
            .I(N__34493));
    LocalMux I__6907 (
            .O(N__34493),
            .I(N__34490));
    Span4Mux_h I__6906 (
            .O(N__34490),
            .I(N__34487));
    Odrv4 I__6905 (
            .O(N__34487),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__6904 (
            .O(N__34484),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__6903 (
            .O(N__34481),
            .I(N__34478));
    LocalMux I__6902 (
            .O(N__34478),
            .I(N__34475));
    Span4Mux_h I__6901 (
            .O(N__34475),
            .I(N__34472));
    Span4Mux_v I__6900 (
            .O(N__34472),
            .I(N__34469));
    Odrv4 I__6899 (
            .O(N__34469),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__6898 (
            .O(N__34466),
            .I(N__34463));
    LocalMux I__6897 (
            .O(N__34463),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__6896 (
            .O(N__34460),
            .I(N__34457));
    LocalMux I__6895 (
            .O(N__34457),
            .I(N__34454));
    Odrv12 I__6894 (
            .O(N__34454),
            .I(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ));
    InMux I__6893 (
            .O(N__34451),
            .I(N__34448));
    LocalMux I__6892 (
            .O(N__34448),
            .I(N__34445));
    Span4Mux_h I__6891 (
            .O(N__34445),
            .I(N__34442));
    Odrv4 I__6890 (
            .O(N__34442),
            .I(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ));
    CascadeMux I__6889 (
            .O(N__34439),
            .I(N__34436));
    InMux I__6888 (
            .O(N__34436),
            .I(N__34433));
    LocalMux I__6887 (
            .O(N__34433),
            .I(N__34430));
    Odrv4 I__6886 (
            .O(N__34430),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__6885 (
            .O(N__34427),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    CascadeMux I__6884 (
            .O(N__34424),
            .I(N__34421));
    InMux I__6883 (
            .O(N__34421),
            .I(N__34418));
    LocalMux I__6882 (
            .O(N__34418),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__6881 (
            .O(N__34415),
            .I(N__34412));
    LocalMux I__6880 (
            .O(N__34412),
            .I(N__34409));
    Odrv4 I__6879 (
            .O(N__34409),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__6878 (
            .O(N__34406),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__6877 (
            .O(N__34403),
            .I(N__34400));
    LocalMux I__6876 (
            .O(N__34400),
            .I(N__34397));
    Odrv4 I__6875 (
            .O(N__34397),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__6874 (
            .O(N__34394),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__6873 (
            .O(N__34391),
            .I(N__34388));
    LocalMux I__6872 (
            .O(N__34388),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__6871 (
            .O(N__34385),
            .I(bfn_14_16_0_));
    InMux I__6870 (
            .O(N__34382),
            .I(N__34379));
    LocalMux I__6869 (
            .O(N__34379),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__6868 (
            .O(N__34376),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__6867 (
            .O(N__34373),
            .I(N__34370));
    LocalMux I__6866 (
            .O(N__34370),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__6865 (
            .O(N__34367),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__6864 (
            .O(N__34364),
            .I(N__34361));
    LocalMux I__6863 (
            .O(N__34361),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__6862 (
            .O(N__34358),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__6861 (
            .O(N__34355),
            .I(N__34352));
    LocalMux I__6860 (
            .O(N__34352),
            .I(N__34349));
    Odrv4 I__6859 (
            .O(N__34349),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__6858 (
            .O(N__34346),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__6857 (
            .O(N__34343),
            .I(N__34340));
    LocalMux I__6856 (
            .O(N__34340),
            .I(N__34337));
    Odrv4 I__6855 (
            .O(N__34337),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__6854 (
            .O(N__34334),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__6853 (
            .O(N__34331),
            .I(N__34328));
    LocalMux I__6852 (
            .O(N__34328),
            .I(N__34325));
    Span4Mux_h I__6851 (
            .O(N__34325),
            .I(N__34322));
    Odrv4 I__6850 (
            .O(N__34322),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__6849 (
            .O(N__34319),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__6848 (
            .O(N__34316),
            .I(N__34313));
    LocalMux I__6847 (
            .O(N__34313),
            .I(N__34310));
    Odrv4 I__6846 (
            .O(N__34310),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    CascadeMux I__6845 (
            .O(N__34307),
            .I(N__34304));
    InMux I__6844 (
            .O(N__34304),
            .I(N__34301));
    LocalMux I__6843 (
            .O(N__34301),
            .I(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ));
    CascadeMux I__6842 (
            .O(N__34298),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_));
    InMux I__6841 (
            .O(N__34295),
            .I(N__34292));
    LocalMux I__6840 (
            .O(N__34292),
            .I(N__34288));
    InMux I__6839 (
            .O(N__34291),
            .I(N__34285));
    Odrv4 I__6838 (
            .O(N__34288),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    LocalMux I__6837 (
            .O(N__34285),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    CascadeMux I__6836 (
            .O(N__34280),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31_cascade_));
    InMux I__6835 (
            .O(N__34277),
            .I(N__34274));
    LocalMux I__6834 (
            .O(N__34274),
            .I(N__34270));
    InMux I__6833 (
            .O(N__34273),
            .I(N__34267));
    Odrv4 I__6832 (
            .O(N__34270),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    LocalMux I__6831 (
            .O(N__34267),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    InMux I__6830 (
            .O(N__34262),
            .I(N__34258));
    InMux I__6829 (
            .O(N__34261),
            .I(N__34255));
    LocalMux I__6828 (
            .O(N__34258),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    LocalMux I__6827 (
            .O(N__34255),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    CascadeMux I__6826 (
            .O(N__34250),
            .I(N__34247));
    InMux I__6825 (
            .O(N__34247),
            .I(N__34244));
    LocalMux I__6824 (
            .O(N__34244),
            .I(N__34241));
    Odrv12 I__6823 (
            .O(N__34241),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__6822 (
            .O(N__34238),
            .I(N__34235));
    InMux I__6821 (
            .O(N__34235),
            .I(N__34232));
    LocalMux I__6820 (
            .O(N__34232),
            .I(N__34229));
    Span4Mux_h I__6819 (
            .O(N__34229),
            .I(N__34226));
    Odrv4 I__6818 (
            .O(N__34226),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__6817 (
            .O(N__34223),
            .I(bfn_14_11_0_));
    InMux I__6816 (
            .O(N__34220),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__6815 (
            .O(N__34217),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__6814 (
            .O(N__34214),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__6813 (
            .O(N__34211),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__6812 (
            .O(N__34208),
            .I(N__34198));
    InMux I__6811 (
            .O(N__34207),
            .I(N__34198));
    InMux I__6810 (
            .O(N__34206),
            .I(N__34198));
    InMux I__6809 (
            .O(N__34205),
            .I(N__34195));
    LocalMux I__6808 (
            .O(N__34198),
            .I(N__34192));
    LocalMux I__6807 (
            .O(N__34195),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__6806 (
            .O(N__34192),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__6805 (
            .O(N__34187),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__6804 (
            .O(N__34184),
            .I(N__34152));
    InMux I__6803 (
            .O(N__34183),
            .I(N__34152));
    InMux I__6802 (
            .O(N__34182),
            .I(N__34152));
    InMux I__6801 (
            .O(N__34181),
            .I(N__34152));
    IoInMux I__6800 (
            .O(N__34180),
            .I(N__34149));
    InMux I__6799 (
            .O(N__34179),
            .I(N__34133));
    InMux I__6798 (
            .O(N__34178),
            .I(N__34133));
    InMux I__6797 (
            .O(N__34177),
            .I(N__34133));
    InMux I__6796 (
            .O(N__34176),
            .I(N__34133));
    InMux I__6795 (
            .O(N__34175),
            .I(N__34126));
    InMux I__6794 (
            .O(N__34174),
            .I(N__34126));
    InMux I__6793 (
            .O(N__34173),
            .I(N__34126));
    InMux I__6792 (
            .O(N__34172),
            .I(N__34117));
    InMux I__6791 (
            .O(N__34171),
            .I(N__34117));
    InMux I__6790 (
            .O(N__34170),
            .I(N__34117));
    InMux I__6789 (
            .O(N__34169),
            .I(N__34117));
    InMux I__6788 (
            .O(N__34168),
            .I(N__34108));
    InMux I__6787 (
            .O(N__34167),
            .I(N__34108));
    InMux I__6786 (
            .O(N__34166),
            .I(N__34108));
    InMux I__6785 (
            .O(N__34165),
            .I(N__34108));
    InMux I__6784 (
            .O(N__34164),
            .I(N__34099));
    InMux I__6783 (
            .O(N__34163),
            .I(N__34099));
    InMux I__6782 (
            .O(N__34162),
            .I(N__34099));
    InMux I__6781 (
            .O(N__34161),
            .I(N__34099));
    LocalMux I__6780 (
            .O(N__34152),
            .I(N__34096));
    LocalMux I__6779 (
            .O(N__34149),
            .I(N__34093));
    InMux I__6778 (
            .O(N__34148),
            .I(N__34083));
    InMux I__6777 (
            .O(N__34147),
            .I(N__34083));
    InMux I__6776 (
            .O(N__34146),
            .I(N__34083));
    InMux I__6775 (
            .O(N__34145),
            .I(N__34083));
    InMux I__6774 (
            .O(N__34144),
            .I(N__34076));
    InMux I__6773 (
            .O(N__34143),
            .I(N__34076));
    InMux I__6772 (
            .O(N__34142),
            .I(N__34076));
    LocalMux I__6771 (
            .O(N__34133),
            .I(N__34073));
    LocalMux I__6770 (
            .O(N__34126),
            .I(N__34064));
    LocalMux I__6769 (
            .O(N__34117),
            .I(N__34064));
    LocalMux I__6768 (
            .O(N__34108),
            .I(N__34064));
    LocalMux I__6767 (
            .O(N__34099),
            .I(N__34064));
    Span4Mux_h I__6766 (
            .O(N__34096),
            .I(N__34061));
    Span4Mux_s0_v I__6765 (
            .O(N__34093),
            .I(N__34058));
    InMux I__6764 (
            .O(N__34092),
            .I(N__34055));
    LocalMux I__6763 (
            .O(N__34083),
            .I(N__34046));
    LocalMux I__6762 (
            .O(N__34076),
            .I(N__34046));
    Span4Mux_v I__6761 (
            .O(N__34073),
            .I(N__34046));
    Span4Mux_v I__6760 (
            .O(N__34064),
            .I(N__34046));
    Span4Mux_v I__6759 (
            .O(N__34061),
            .I(N__34041));
    Span4Mux_v I__6758 (
            .O(N__34058),
            .I(N__34041));
    LocalMux I__6757 (
            .O(N__34055),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__6756 (
            .O(N__34046),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    Odrv4 I__6755 (
            .O(N__34041),
            .I(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ));
    InMux I__6754 (
            .O(N__34034),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    CascadeMux I__6753 (
            .O(N__34031),
            .I(N__34027));
    CascadeMux I__6752 (
            .O(N__34030),
            .I(N__34024));
    InMux I__6751 (
            .O(N__34027),
            .I(N__34016));
    InMux I__6750 (
            .O(N__34024),
            .I(N__34016));
    InMux I__6749 (
            .O(N__34023),
            .I(N__34016));
    LocalMux I__6748 (
            .O(N__34016),
            .I(N__34012));
    InMux I__6747 (
            .O(N__34015),
            .I(N__34009));
    Span4Mux_v I__6746 (
            .O(N__34012),
            .I(N__34006));
    LocalMux I__6745 (
            .O(N__34009),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__6744 (
            .O(N__34006),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__6743 (
            .O(N__34001),
            .I(N__33998));
    LocalMux I__6742 (
            .O(N__33998),
            .I(N__33994));
    InMux I__6741 (
            .O(N__33997),
            .I(N__33991));
    Odrv4 I__6740 (
            .O(N__33994),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    LocalMux I__6739 (
            .O(N__33991),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    InMux I__6738 (
            .O(N__33986),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__6737 (
            .O(N__33983),
            .I(bfn_14_10_0_));
    InMux I__6736 (
            .O(N__33980),
            .I(N__33973));
    InMux I__6735 (
            .O(N__33979),
            .I(N__33973));
    InMux I__6734 (
            .O(N__33978),
            .I(N__33970));
    LocalMux I__6733 (
            .O(N__33973),
            .I(N__33967));
    LocalMux I__6732 (
            .O(N__33970),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__6731 (
            .O(N__33967),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__6730 (
            .O(N__33962),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    CascadeMux I__6729 (
            .O(N__33959),
            .I(N__33956));
    InMux I__6728 (
            .O(N__33956),
            .I(N__33949));
    InMux I__6727 (
            .O(N__33955),
            .I(N__33949));
    InMux I__6726 (
            .O(N__33954),
            .I(N__33946));
    LocalMux I__6725 (
            .O(N__33949),
            .I(N__33943));
    LocalMux I__6724 (
            .O(N__33946),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__6723 (
            .O(N__33943),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__6722 (
            .O(N__33938),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__6721 (
            .O(N__33935),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__6720 (
            .O(N__33932),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__6719 (
            .O(N__33929),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__6718 (
            .O(N__33926),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    InMux I__6717 (
            .O(N__33923),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__6716 (
            .O(N__33920),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__6715 (
            .O(N__33917),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__6714 (
            .O(N__33914),
            .I(bfn_14_9_0_));
    InMux I__6713 (
            .O(N__33911),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__6712 (
            .O(N__33908),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__6711 (
            .O(N__33905),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__6710 (
            .O(N__33902),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__6709 (
            .O(N__33899),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__6708 (
            .O(N__33896),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    CascadeMux I__6707 (
            .O(N__33893),
            .I(N__33890));
    InMux I__6706 (
            .O(N__33890),
            .I(N__33884));
    InMux I__6705 (
            .O(N__33889),
            .I(N__33884));
    LocalMux I__6704 (
            .O(N__33884),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__6703 (
            .O(N__33881),
            .I(N__33878));
    LocalMux I__6702 (
            .O(N__33878),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ));
    InMux I__6701 (
            .O(N__33875),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__6700 (
            .O(N__33872),
            .I(N__33869));
    InMux I__6699 (
            .O(N__33869),
            .I(N__33866));
    LocalMux I__6698 (
            .O(N__33866),
            .I(N__33863));
    Odrv4 I__6697 (
            .O(N__33863),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ));
    InMux I__6696 (
            .O(N__33860),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__6695 (
            .O(N__33857),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__6694 (
            .O(N__33854),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__6693 (
            .O(N__33851),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__6692 (
            .O(N__33848),
            .I(N__33842));
    InMux I__6691 (
            .O(N__33847),
            .I(N__33842));
    LocalMux I__6690 (
            .O(N__33842),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    InMux I__6689 (
            .O(N__33839),
            .I(N__33836));
    LocalMux I__6688 (
            .O(N__33836),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__6687 (
            .O(N__33833),
            .I(N__33830));
    LocalMux I__6686 (
            .O(N__33830),
            .I(N__33827));
    Span4Mux_h I__6685 (
            .O(N__33827),
            .I(N__33824));
    Odrv4 I__6684 (
            .O(N__33824),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__6683 (
            .O(N__33821),
            .I(N__33818));
    LocalMux I__6682 (
            .O(N__33818),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__6681 (
            .O(N__33815),
            .I(N__33812));
    LocalMux I__6680 (
            .O(N__33812),
            .I(N__33809));
    Span4Mux_v I__6679 (
            .O(N__33809),
            .I(N__33806));
    Odrv4 I__6678 (
            .O(N__33806),
            .I(\current_shift_inst.control_input_axb_10 ));
    CascadeMux I__6677 (
            .O(N__33803),
            .I(N__33800));
    InMux I__6676 (
            .O(N__33800),
            .I(N__33797));
    LocalMux I__6675 (
            .O(N__33797),
            .I(N__33794));
    Odrv4 I__6674 (
            .O(N__33794),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__6673 (
            .O(N__33791),
            .I(N__33788));
    LocalMux I__6672 (
            .O(N__33788),
            .I(N__33784));
    InMux I__6671 (
            .O(N__33787),
            .I(N__33781));
    Span4Mux_v I__6670 (
            .O(N__33784),
            .I(N__33778));
    LocalMux I__6669 (
            .O(N__33781),
            .I(N__33775));
    Span4Mux_v I__6668 (
            .O(N__33778),
            .I(N__33772));
    Span4Mux_v I__6667 (
            .O(N__33775),
            .I(N__33769));
    Odrv4 I__6666 (
            .O(N__33772),
            .I(state_ns_i_a2_1));
    Odrv4 I__6665 (
            .O(N__33769),
            .I(state_ns_i_a2_1));
    InMux I__6664 (
            .O(N__33764),
            .I(N__33757));
    InMux I__6663 (
            .O(N__33763),
            .I(N__33757));
    InMux I__6662 (
            .O(N__33762),
            .I(N__33754));
    LocalMux I__6661 (
            .O(N__33757),
            .I(N__33751));
    LocalMux I__6660 (
            .O(N__33754),
            .I(N__33748));
    Span4Mux_v I__6659 (
            .O(N__33751),
            .I(N__33745));
    Span4Mux_h I__6658 (
            .O(N__33748),
            .I(N__33742));
    Sp12to4 I__6657 (
            .O(N__33745),
            .I(N__33738));
    Span4Mux_h I__6656 (
            .O(N__33742),
            .I(N__33735));
    InMux I__6655 (
            .O(N__33741),
            .I(N__33732));
    Span12Mux_h I__6654 (
            .O(N__33738),
            .I(N__33729));
    Odrv4 I__6653 (
            .O(N__33735),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__6652 (
            .O(N__33732),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv12 I__6651 (
            .O(N__33729),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__6650 (
            .O(N__33722),
            .I(N__33719));
    LocalMux I__6649 (
            .O(N__33719),
            .I(\phase_controller_inst1.start_timer_hc_0_sqmuxa ));
    CascadeMux I__6648 (
            .O(N__33716),
            .I(N__33712));
    InMux I__6647 (
            .O(N__33715),
            .I(N__33709));
    InMux I__6646 (
            .O(N__33712),
            .I(N__33705));
    LocalMux I__6645 (
            .O(N__33709),
            .I(N__33702));
    InMux I__6644 (
            .O(N__33708),
            .I(N__33699));
    LocalMux I__6643 (
            .O(N__33705),
            .I(N__33692));
    Span4Mux_v I__6642 (
            .O(N__33702),
            .I(N__33692));
    LocalMux I__6641 (
            .O(N__33699),
            .I(N__33692));
    Span4Mux_v I__6640 (
            .O(N__33692),
            .I(N__33689));
    Odrv4 I__6639 (
            .O(N__33689),
            .I(il_max_comp1_D2));
    IoInMux I__6638 (
            .O(N__33686),
            .I(N__33683));
    LocalMux I__6637 (
            .O(N__33683),
            .I(N__33680));
    Odrv12 I__6636 (
            .O(N__33680),
            .I(\current_shift_inst.timer_s1.N_162_i ));
    InMux I__6635 (
            .O(N__33677),
            .I(N__33674));
    LocalMux I__6634 (
            .O(N__33674),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__6633 (
            .O(N__33671),
            .I(N__33668));
    LocalMux I__6632 (
            .O(N__33668),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__6631 (
            .O(N__33665),
            .I(N__33662));
    LocalMux I__6630 (
            .O(N__33662),
            .I(N__33659));
    Span4Mux_v I__6629 (
            .O(N__33659),
            .I(N__33656));
    Odrv4 I__6628 (
            .O(N__33656),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__6627 (
            .O(N__33653),
            .I(N__33650));
    LocalMux I__6626 (
            .O(N__33650),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__6625 (
            .O(N__33647),
            .I(N__33644));
    LocalMux I__6624 (
            .O(N__33644),
            .I(N__33641));
    Span4Mux_v I__6623 (
            .O(N__33641),
            .I(N__33638));
    Odrv4 I__6622 (
            .O(N__33638),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__6621 (
            .O(N__33635),
            .I(N__33632));
    LocalMux I__6620 (
            .O(N__33632),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__6619 (
            .O(N__33629),
            .I(N__33626));
    LocalMux I__6618 (
            .O(N__33626),
            .I(N__33623));
    Span4Mux_h I__6617 (
            .O(N__33623),
            .I(N__33620));
    Odrv4 I__6616 (
            .O(N__33620),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__6615 (
            .O(N__33617),
            .I(N__33614));
    LocalMux I__6614 (
            .O(N__33614),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__6613 (
            .O(N__33611),
            .I(N__33608));
    LocalMux I__6612 (
            .O(N__33608),
            .I(N__33605));
    Span4Mux_h I__6611 (
            .O(N__33605),
            .I(N__33602));
    Odrv4 I__6610 (
            .O(N__33602),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__6609 (
            .O(N__33599),
            .I(N__33596));
    LocalMux I__6608 (
            .O(N__33596),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__6607 (
            .O(N__33593),
            .I(N__33590));
    LocalMux I__6606 (
            .O(N__33590),
            .I(N__33587));
    Span4Mux_h I__6605 (
            .O(N__33587),
            .I(N__33584));
    Odrv4 I__6604 (
            .O(N__33584),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__6603 (
            .O(N__33581),
            .I(N__33578));
    LocalMux I__6602 (
            .O(N__33578),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__6601 (
            .O(N__33575),
            .I(N__33572));
    LocalMux I__6600 (
            .O(N__33572),
            .I(N__33569));
    Span4Mux_h I__6599 (
            .O(N__33569),
            .I(N__33566));
    Odrv4 I__6598 (
            .O(N__33566),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__6597 (
            .O(N__33563),
            .I(N__33560));
    LocalMux I__6596 (
            .O(N__33560),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__6595 (
            .O(N__33557),
            .I(N__33554));
    LocalMux I__6594 (
            .O(N__33554),
            .I(N__33551));
    Span4Mux_h I__6593 (
            .O(N__33551),
            .I(N__33548));
    Odrv4 I__6592 (
            .O(N__33548),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__6591 (
            .O(N__33545),
            .I(N__33542));
    LocalMux I__6590 (
            .O(N__33542),
            .I(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ));
    CascadeMux I__6589 (
            .O(N__33539),
            .I(N__33536));
    InMux I__6588 (
            .O(N__33536),
            .I(N__33533));
    LocalMux I__6587 (
            .O(N__33533),
            .I(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ));
    CascadeMux I__6586 (
            .O(N__33530),
            .I(N__33527));
    InMux I__6585 (
            .O(N__33527),
            .I(N__33524));
    LocalMux I__6584 (
            .O(N__33524),
            .I(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ));
    InMux I__6583 (
            .O(N__33521),
            .I(N__33518));
    LocalMux I__6582 (
            .O(N__33518),
            .I(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ));
    CascadeMux I__6581 (
            .O(N__33515),
            .I(N__33512));
    InMux I__6580 (
            .O(N__33512),
            .I(N__33509));
    LocalMux I__6579 (
            .O(N__33509),
            .I(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ));
    CascadeMux I__6578 (
            .O(N__33506),
            .I(N__33503));
    InMux I__6577 (
            .O(N__33503),
            .I(N__33500));
    LocalMux I__6576 (
            .O(N__33500),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__6575 (
            .O(N__33497),
            .I(N__33494));
    LocalMux I__6574 (
            .O(N__33494),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__6573 (
            .O(N__33491),
            .I(N__33488));
    LocalMux I__6572 (
            .O(N__33488),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__6571 (
            .O(N__33485),
            .I(N__33482));
    LocalMux I__6570 (
            .O(N__33482),
            .I(N__33479));
    Span4Mux_h I__6569 (
            .O(N__33479),
            .I(N__33476));
    Odrv4 I__6568 (
            .O(N__33476),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__6567 (
            .O(N__33473),
            .I(N__33470));
    LocalMux I__6566 (
            .O(N__33470),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    CascadeMux I__6565 (
            .O(N__33467),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ));
    CascadeMux I__6564 (
            .O(N__33464),
            .I(N__33460));
    InMux I__6563 (
            .O(N__33463),
            .I(N__33457));
    InMux I__6562 (
            .O(N__33460),
            .I(N__33454));
    LocalMux I__6561 (
            .O(N__33457),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    LocalMux I__6560 (
            .O(N__33454),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    InMux I__6559 (
            .O(N__33449),
            .I(N__33446));
    LocalMux I__6558 (
            .O(N__33446),
            .I(N__33440));
    InMux I__6557 (
            .O(N__33445),
            .I(N__33437));
    InMux I__6556 (
            .O(N__33444),
            .I(N__33432));
    InMux I__6555 (
            .O(N__33443),
            .I(N__33432));
    Span4Mux_h I__6554 (
            .O(N__33440),
            .I(N__33429));
    LocalMux I__6553 (
            .O(N__33437),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__6552 (
            .O(N__33432),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__6551 (
            .O(N__33429),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__6550 (
            .O(N__33422),
            .I(N__33384));
    InMux I__6549 (
            .O(N__33421),
            .I(N__33384));
    InMux I__6548 (
            .O(N__33420),
            .I(N__33384));
    InMux I__6547 (
            .O(N__33419),
            .I(N__33384));
    InMux I__6546 (
            .O(N__33418),
            .I(N__33375));
    InMux I__6545 (
            .O(N__33417),
            .I(N__33375));
    InMux I__6544 (
            .O(N__33416),
            .I(N__33375));
    InMux I__6543 (
            .O(N__33415),
            .I(N__33375));
    InMux I__6542 (
            .O(N__33414),
            .I(N__33370));
    InMux I__6541 (
            .O(N__33413),
            .I(N__33370));
    InMux I__6540 (
            .O(N__33412),
            .I(N__33361));
    InMux I__6539 (
            .O(N__33411),
            .I(N__33361));
    InMux I__6538 (
            .O(N__33410),
            .I(N__33361));
    InMux I__6537 (
            .O(N__33409),
            .I(N__33361));
    InMux I__6536 (
            .O(N__33408),
            .I(N__33352));
    InMux I__6535 (
            .O(N__33407),
            .I(N__33352));
    InMux I__6534 (
            .O(N__33406),
            .I(N__33352));
    InMux I__6533 (
            .O(N__33405),
            .I(N__33352));
    InMux I__6532 (
            .O(N__33404),
            .I(N__33343));
    InMux I__6531 (
            .O(N__33403),
            .I(N__33343));
    InMux I__6530 (
            .O(N__33402),
            .I(N__33343));
    InMux I__6529 (
            .O(N__33401),
            .I(N__33343));
    InMux I__6528 (
            .O(N__33400),
            .I(N__33334));
    InMux I__6527 (
            .O(N__33399),
            .I(N__33334));
    InMux I__6526 (
            .O(N__33398),
            .I(N__33334));
    InMux I__6525 (
            .O(N__33397),
            .I(N__33334));
    InMux I__6524 (
            .O(N__33396),
            .I(N__33325));
    InMux I__6523 (
            .O(N__33395),
            .I(N__33325));
    InMux I__6522 (
            .O(N__33394),
            .I(N__33325));
    InMux I__6521 (
            .O(N__33393),
            .I(N__33325));
    LocalMux I__6520 (
            .O(N__33384),
            .I(N__33322));
    LocalMux I__6519 (
            .O(N__33375),
            .I(N__33319));
    LocalMux I__6518 (
            .O(N__33370),
            .I(N__33314));
    LocalMux I__6517 (
            .O(N__33361),
            .I(N__33314));
    LocalMux I__6516 (
            .O(N__33352),
            .I(N__33305));
    LocalMux I__6515 (
            .O(N__33343),
            .I(N__33305));
    LocalMux I__6514 (
            .O(N__33334),
            .I(N__33305));
    LocalMux I__6513 (
            .O(N__33325),
            .I(N__33305));
    Odrv4 I__6512 (
            .O(N__33322),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__6511 (
            .O(N__33319),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__6510 (
            .O(N__33314),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv12 I__6509 (
            .O(N__33305),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__6508 (
            .O(N__33296),
            .I(N__33293));
    LocalMux I__6507 (
            .O(N__33293),
            .I(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ));
    CascadeMux I__6506 (
            .O(N__33290),
            .I(N__33287));
    InMux I__6505 (
            .O(N__33287),
            .I(N__33284));
    LocalMux I__6504 (
            .O(N__33284),
            .I(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ));
    InMux I__6503 (
            .O(N__33281),
            .I(N__33278));
    LocalMux I__6502 (
            .O(N__33278),
            .I(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ));
    InMux I__6501 (
            .O(N__33275),
            .I(N__33272));
    LocalMux I__6500 (
            .O(N__33272),
            .I(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ));
    CascadeMux I__6499 (
            .O(N__33269),
            .I(N__33266));
    InMux I__6498 (
            .O(N__33266),
            .I(N__33263));
    LocalMux I__6497 (
            .O(N__33263),
            .I(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ));
    InMux I__6496 (
            .O(N__33260),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__6495 (
            .O(N__33257),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__6494 (
            .O(N__33254),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__6493 (
            .O(N__33251),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__6492 (
            .O(N__33248),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    CEMux I__6491 (
            .O(N__33245),
            .I(N__33241));
    CEMux I__6490 (
            .O(N__33244),
            .I(N__33238));
    LocalMux I__6489 (
            .O(N__33241),
            .I(N__33233));
    LocalMux I__6488 (
            .O(N__33238),
            .I(N__33230));
    CEMux I__6487 (
            .O(N__33237),
            .I(N__33227));
    CEMux I__6486 (
            .O(N__33236),
            .I(N__33224));
    Span4Mux_v I__6485 (
            .O(N__33233),
            .I(N__33217));
    Span4Mux_h I__6484 (
            .O(N__33230),
            .I(N__33217));
    LocalMux I__6483 (
            .O(N__33227),
            .I(N__33217));
    LocalMux I__6482 (
            .O(N__33224),
            .I(N__33214));
    Span4Mux_v I__6481 (
            .O(N__33217),
            .I(N__33211));
    Span4Mux_h I__6480 (
            .O(N__33214),
            .I(N__33208));
    Odrv4 I__6479 (
            .O(N__33211),
            .I(\delay_measurement_inst.delay_tr_timer.N_205_i ));
    Odrv4 I__6478 (
            .O(N__33208),
            .I(\delay_measurement_inst.delay_tr_timer.N_205_i ));
    CascadeMux I__6477 (
            .O(N__33203),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    CascadeMux I__6476 (
            .O(N__33200),
            .I(N__33196));
    InMux I__6475 (
            .O(N__33199),
            .I(N__33191));
    InMux I__6474 (
            .O(N__33196),
            .I(N__33184));
    InMux I__6473 (
            .O(N__33195),
            .I(N__33184));
    InMux I__6472 (
            .O(N__33194),
            .I(N__33184));
    LocalMux I__6471 (
            .O(N__33191),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6470 (
            .O(N__33184),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    InMux I__6469 (
            .O(N__33179),
            .I(N__33176));
    LocalMux I__6468 (
            .O(N__33176),
            .I(\current_shift_inst.un4_control_input1_1 ));
    InMux I__6467 (
            .O(N__33173),
            .I(bfn_13_12_0_));
    InMux I__6466 (
            .O(N__33170),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__6465 (
            .O(N__33167),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__6464 (
            .O(N__33164),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__6463 (
            .O(N__33161),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__6462 (
            .O(N__33158),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__6461 (
            .O(N__33155),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__6460 (
            .O(N__33152),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__6459 (
            .O(N__33149),
            .I(bfn_13_13_0_));
    InMux I__6458 (
            .O(N__33146),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__6457 (
            .O(N__33143),
            .I(bfn_13_11_0_));
    InMux I__6456 (
            .O(N__33140),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__6455 (
            .O(N__33137),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__6454 (
            .O(N__33134),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__6453 (
            .O(N__33131),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__6452 (
            .O(N__33128),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__6451 (
            .O(N__33125),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__6450 (
            .O(N__33122),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    CascadeMux I__6449 (
            .O(N__33119),
            .I(N__33115));
    InMux I__6448 (
            .O(N__33118),
            .I(N__33107));
    InMux I__6447 (
            .O(N__33115),
            .I(N__33107));
    InMux I__6446 (
            .O(N__33114),
            .I(N__33107));
    LocalMux I__6445 (
            .O(N__33107),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    InMux I__6444 (
            .O(N__33104),
            .I(bfn_13_10_0_));
    InMux I__6443 (
            .O(N__33101),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__6442 (
            .O(N__33098),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__6441 (
            .O(N__33095),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__6440 (
            .O(N__33092),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__6439 (
            .O(N__33089),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__6438 (
            .O(N__33086),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__6437 (
            .O(N__33083),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ));
    InMux I__6436 (
            .O(N__33080),
            .I(N__33073));
    InMux I__6435 (
            .O(N__33079),
            .I(N__33068));
    InMux I__6434 (
            .O(N__33078),
            .I(N__33068));
    InMux I__6433 (
            .O(N__33077),
            .I(N__33065));
    InMux I__6432 (
            .O(N__33076),
            .I(N__33062));
    LocalMux I__6431 (
            .O(N__33073),
            .I(N__33057));
    LocalMux I__6430 (
            .O(N__33068),
            .I(N__33057));
    LocalMux I__6429 (
            .O(N__33065),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    LocalMux I__6428 (
            .O(N__33062),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    Odrv4 I__6427 (
            .O(N__33057),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__6426 (
            .O(N__33050),
            .I(N__33046));
    InMux I__6425 (
            .O(N__33049),
            .I(N__33043));
    LocalMux I__6424 (
            .O(N__33046),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    LocalMux I__6423 (
            .O(N__33043),
            .I(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ));
    CascadeMux I__6422 (
            .O(N__33038),
            .I(N__33035));
    InMux I__6421 (
            .O(N__33035),
            .I(N__33032));
    LocalMux I__6420 (
            .O(N__33032),
            .I(N__33029));
    Odrv4 I__6419 (
            .O(N__33029),
            .I(\phase_controller_inst2.stoper_tr.un4_running_df30 ));
    InMux I__6418 (
            .O(N__33026),
            .I(N__33017));
    InMux I__6417 (
            .O(N__33025),
            .I(N__33017));
    InMux I__6416 (
            .O(N__33024),
            .I(N__33017));
    LocalMux I__6415 (
            .O(N__33017),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    CascadeMux I__6414 (
            .O(N__33014),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_));
    InMux I__6413 (
            .O(N__33011),
            .I(N__33007));
    CascadeMux I__6412 (
            .O(N__33010),
            .I(N__33004));
    LocalMux I__6411 (
            .O(N__33007),
            .I(N__32999));
    InMux I__6410 (
            .O(N__33004),
            .I(N__32996));
    InMux I__6409 (
            .O(N__33003),
            .I(N__32991));
    InMux I__6408 (
            .O(N__33002),
            .I(N__32991));
    Span12Mux_v I__6407 (
            .O(N__32999),
            .I(N__32988));
    LocalMux I__6406 (
            .O(N__32996),
            .I(N__32985));
    LocalMux I__6405 (
            .O(N__32991),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv12 I__6404 (
            .O(N__32988),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__6403 (
            .O(N__32985),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    IoInMux I__6402 (
            .O(N__32978),
            .I(N__32975));
    LocalMux I__6401 (
            .O(N__32975),
            .I(N__32972));
    IoSpan4Mux I__6400 (
            .O(N__32972),
            .I(N__32969));
    Sp12to4 I__6399 (
            .O(N__32969),
            .I(N__32966));
    Odrv12 I__6398 (
            .O(N__32966),
            .I(s4_phy_c));
    InMux I__6397 (
            .O(N__32963),
            .I(N__32960));
    LocalMux I__6396 (
            .O(N__32960),
            .I(N__32956));
    InMux I__6395 (
            .O(N__32959),
            .I(N__32953));
    Span4Mux_h I__6394 (
            .O(N__32956),
            .I(N__32948));
    LocalMux I__6393 (
            .O(N__32953),
            .I(N__32948));
    Span4Mux_h I__6392 (
            .O(N__32948),
            .I(N__32943));
    InMux I__6391 (
            .O(N__32947),
            .I(N__32940));
    InMux I__6390 (
            .O(N__32946),
            .I(N__32937));
    Span4Mux_v I__6389 (
            .O(N__32943),
            .I(N__32934));
    LocalMux I__6388 (
            .O(N__32940),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    LocalMux I__6387 (
            .O(N__32937),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__6386 (
            .O(N__32934),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    ClkMux I__6385 (
            .O(N__32927),
            .I(N__32921));
    ClkMux I__6384 (
            .O(N__32926),
            .I(N__32921));
    GlobalMux I__6383 (
            .O(N__32921),
            .I(N__32918));
    gio2CtrlBuf I__6382 (
            .O(N__32918),
            .I(delay_hc_input_c_g));
    IoInMux I__6381 (
            .O(N__32915),
            .I(N__32912));
    LocalMux I__6380 (
            .O(N__32912),
            .I(N__32909));
    Span4Mux_s0_v I__6379 (
            .O(N__32909),
            .I(N__32906));
    Odrv4 I__6378 (
            .O(N__32906),
            .I(\pll_inst.red_c_i ));
    InMux I__6377 (
            .O(N__32903),
            .I(N__32899));
    InMux I__6376 (
            .O(N__32902),
            .I(N__32896));
    LocalMux I__6375 (
            .O(N__32899),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__6374 (
            .O(N__32896),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__6373 (
            .O(N__32891),
            .I(N__32887));
    InMux I__6372 (
            .O(N__32890),
            .I(N__32884));
    LocalMux I__6371 (
            .O(N__32887),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    LocalMux I__6370 (
            .O(N__32884),
            .I(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ));
    InMux I__6369 (
            .O(N__32879),
            .I(N__32875));
    CascadeMux I__6368 (
            .O(N__32878),
            .I(N__32872));
    LocalMux I__6367 (
            .O(N__32875),
            .I(N__32867));
    InMux I__6366 (
            .O(N__32872),
            .I(N__32864));
    InMux I__6365 (
            .O(N__32871),
            .I(N__32859));
    InMux I__6364 (
            .O(N__32870),
            .I(N__32859));
    Odrv4 I__6363 (
            .O(N__32867),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__6362 (
            .O(N__32864),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__6361 (
            .O(N__32859),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    CascadeMux I__6360 (
            .O(N__32852),
            .I(N__32848));
    InMux I__6359 (
            .O(N__32851),
            .I(N__32844));
    InMux I__6358 (
            .O(N__32848),
            .I(N__32841));
    InMux I__6357 (
            .O(N__32847),
            .I(N__32838));
    LocalMux I__6356 (
            .O(N__32844),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__6355 (
            .O(N__32841),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__6354 (
            .O(N__32838),
            .I(\phase_controller_inst2.tr_time_passed ));
    CascadeMux I__6353 (
            .O(N__32831),
            .I(N__32827));
    InMux I__6352 (
            .O(N__32830),
            .I(N__32824));
    InMux I__6351 (
            .O(N__32827),
            .I(N__32821));
    LocalMux I__6350 (
            .O(N__32824),
            .I(N__32818));
    LocalMux I__6349 (
            .O(N__32821),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    Odrv4 I__6348 (
            .O(N__32818),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    CascadeMux I__6347 (
            .O(N__32813),
            .I(N__32808));
    InMux I__6346 (
            .O(N__32812),
            .I(N__32803));
    InMux I__6345 (
            .O(N__32811),
            .I(N__32803));
    InMux I__6344 (
            .O(N__32808),
            .I(N__32798));
    LocalMux I__6343 (
            .O(N__32803),
            .I(N__32795));
    InMux I__6342 (
            .O(N__32802),
            .I(N__32790));
    InMux I__6341 (
            .O(N__32801),
            .I(N__32790));
    LocalMux I__6340 (
            .O(N__32798),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__6339 (
            .O(N__32795),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    LocalMux I__6338 (
            .O(N__32790),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__6337 (
            .O(N__32783),
            .I(N__32780));
    LocalMux I__6336 (
            .O(N__32780),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__6335 (
            .O(N__32777),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__6334 (
            .O(N__32774),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__6333 (
            .O(N__32771),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__6332 (
            .O(N__32768),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__6331 (
            .O(N__32765),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__6330 (
            .O(N__32762),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__6329 (
            .O(N__32759),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__6328 (
            .O(N__32756),
            .I(N__32753));
    LocalMux I__6327 (
            .O(N__32753),
            .I(N__32750));
    Span4Mux_v I__6326 (
            .O(N__32750),
            .I(N__32747));
    Span4Mux_h I__6325 (
            .O(N__32747),
            .I(N__32744));
    Sp12to4 I__6324 (
            .O(N__32744),
            .I(N__32741));
    Span12Mux_v I__6323 (
            .O(N__32741),
            .I(N__32738));
    Odrv12 I__6322 (
            .O(N__32738),
            .I(il_min_comp1_c));
    InMux I__6321 (
            .O(N__32735),
            .I(N__32732));
    LocalMux I__6320 (
            .O(N__32732),
            .I(il_min_comp1_D1));
    InMux I__6319 (
            .O(N__32729),
            .I(N__32726));
    LocalMux I__6318 (
            .O(N__32726),
            .I(N__32723));
    Odrv4 I__6317 (
            .O(N__32723),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__6316 (
            .O(N__32720),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__6315 (
            .O(N__32717),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    CascadeMux I__6314 (
            .O(N__32714),
            .I(N__32711));
    InMux I__6313 (
            .O(N__32711),
            .I(N__32708));
    LocalMux I__6312 (
            .O(N__32708),
            .I(N__32705));
    Odrv4 I__6311 (
            .O(N__32705),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__6310 (
            .O(N__32702),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__6309 (
            .O(N__32699),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__6308 (
            .O(N__32696),
            .I(bfn_12_18_0_));
    CascadeMux I__6307 (
            .O(N__32693),
            .I(N__32690));
    InMux I__6306 (
            .O(N__32690),
            .I(N__32687));
    LocalMux I__6305 (
            .O(N__32687),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__6304 (
            .O(N__32684),
            .I(N__32681));
    LocalMux I__6303 (
            .O(N__32681),
            .I(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ));
    InMux I__6302 (
            .O(N__32678),
            .I(N__32675));
    LocalMux I__6301 (
            .O(N__32675),
            .I(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ));
    CEMux I__6300 (
            .O(N__32672),
            .I(N__32649));
    CEMux I__6299 (
            .O(N__32671),
            .I(N__32644));
    InMux I__6298 (
            .O(N__32670),
            .I(N__32635));
    InMux I__6297 (
            .O(N__32669),
            .I(N__32635));
    InMux I__6296 (
            .O(N__32668),
            .I(N__32635));
    InMux I__6295 (
            .O(N__32667),
            .I(N__32635));
    InMux I__6294 (
            .O(N__32666),
            .I(N__32626));
    InMux I__6293 (
            .O(N__32665),
            .I(N__32626));
    InMux I__6292 (
            .O(N__32664),
            .I(N__32626));
    InMux I__6291 (
            .O(N__32663),
            .I(N__32626));
    InMux I__6290 (
            .O(N__32662),
            .I(N__32617));
    InMux I__6289 (
            .O(N__32661),
            .I(N__32617));
    InMux I__6288 (
            .O(N__32660),
            .I(N__32617));
    InMux I__6287 (
            .O(N__32659),
            .I(N__32617));
    CEMux I__6286 (
            .O(N__32658),
            .I(N__32613));
    CEMux I__6285 (
            .O(N__32657),
            .I(N__32602));
    CEMux I__6284 (
            .O(N__32656),
            .I(N__32595));
    CEMux I__6283 (
            .O(N__32655),
            .I(N__32591));
    CEMux I__6282 (
            .O(N__32654),
            .I(N__32587));
    CEMux I__6281 (
            .O(N__32653),
            .I(N__32584));
    CEMux I__6280 (
            .O(N__32652),
            .I(N__32581));
    LocalMux I__6279 (
            .O(N__32649),
            .I(N__32578));
    CEMux I__6278 (
            .O(N__32648),
            .I(N__32575));
    CEMux I__6277 (
            .O(N__32647),
            .I(N__32568));
    LocalMux I__6276 (
            .O(N__32644),
            .I(N__32559));
    LocalMux I__6275 (
            .O(N__32635),
            .I(N__32559));
    LocalMux I__6274 (
            .O(N__32626),
            .I(N__32559));
    LocalMux I__6273 (
            .O(N__32617),
            .I(N__32559));
    CEMux I__6272 (
            .O(N__32616),
            .I(N__32556));
    LocalMux I__6271 (
            .O(N__32613),
            .I(N__32549));
    InMux I__6270 (
            .O(N__32612),
            .I(N__32540));
    InMux I__6269 (
            .O(N__32611),
            .I(N__32540));
    InMux I__6268 (
            .O(N__32610),
            .I(N__32540));
    InMux I__6267 (
            .O(N__32609),
            .I(N__32540));
    InMux I__6266 (
            .O(N__32608),
            .I(N__32531));
    InMux I__6265 (
            .O(N__32607),
            .I(N__32531));
    InMux I__6264 (
            .O(N__32606),
            .I(N__32531));
    InMux I__6263 (
            .O(N__32605),
            .I(N__32531));
    LocalMux I__6262 (
            .O(N__32602),
            .I(N__32528));
    CEMux I__6261 (
            .O(N__32601),
            .I(N__32525));
    InMux I__6260 (
            .O(N__32600),
            .I(N__32518));
    InMux I__6259 (
            .O(N__32599),
            .I(N__32518));
    InMux I__6258 (
            .O(N__32598),
            .I(N__32518));
    LocalMux I__6257 (
            .O(N__32595),
            .I(N__32515));
    CEMux I__6256 (
            .O(N__32594),
            .I(N__32512));
    LocalMux I__6255 (
            .O(N__32591),
            .I(N__32509));
    CEMux I__6254 (
            .O(N__32590),
            .I(N__32506));
    LocalMux I__6253 (
            .O(N__32587),
            .I(N__32503));
    LocalMux I__6252 (
            .O(N__32584),
            .I(N__32498));
    LocalMux I__6251 (
            .O(N__32581),
            .I(N__32498));
    Span4Mux_s3_v I__6250 (
            .O(N__32578),
            .I(N__32492));
    LocalMux I__6249 (
            .O(N__32575),
            .I(N__32492));
    CEMux I__6248 (
            .O(N__32574),
            .I(N__32489));
    InMux I__6247 (
            .O(N__32573),
            .I(N__32482));
    InMux I__6246 (
            .O(N__32572),
            .I(N__32482));
    InMux I__6245 (
            .O(N__32571),
            .I(N__32482));
    LocalMux I__6244 (
            .O(N__32568),
            .I(N__32475));
    Span4Mux_v I__6243 (
            .O(N__32559),
            .I(N__32475));
    LocalMux I__6242 (
            .O(N__32556),
            .I(N__32475));
    InMux I__6241 (
            .O(N__32555),
            .I(N__32466));
    InMux I__6240 (
            .O(N__32554),
            .I(N__32466));
    InMux I__6239 (
            .O(N__32553),
            .I(N__32466));
    InMux I__6238 (
            .O(N__32552),
            .I(N__32466));
    Span4Mux_h I__6237 (
            .O(N__32549),
            .I(N__32453));
    LocalMux I__6236 (
            .O(N__32540),
            .I(N__32453));
    LocalMux I__6235 (
            .O(N__32531),
            .I(N__32453));
    Span4Mux_s3_v I__6234 (
            .O(N__32528),
            .I(N__32453));
    LocalMux I__6233 (
            .O(N__32525),
            .I(N__32453));
    LocalMux I__6232 (
            .O(N__32518),
            .I(N__32453));
    Span4Mux_v I__6231 (
            .O(N__32515),
            .I(N__32448));
    LocalMux I__6230 (
            .O(N__32512),
            .I(N__32448));
    Span4Mux_v I__6229 (
            .O(N__32509),
            .I(N__32443));
    LocalMux I__6228 (
            .O(N__32506),
            .I(N__32443));
    Span4Mux_v I__6227 (
            .O(N__32503),
            .I(N__32438));
    Span4Mux_v I__6226 (
            .O(N__32498),
            .I(N__32438));
    InMux I__6225 (
            .O(N__32497),
            .I(N__32435));
    Span4Mux_v I__6224 (
            .O(N__32492),
            .I(N__32432));
    LocalMux I__6223 (
            .O(N__32489),
            .I(N__32419));
    LocalMux I__6222 (
            .O(N__32482),
            .I(N__32419));
    Span4Mux_v I__6221 (
            .O(N__32475),
            .I(N__32419));
    LocalMux I__6220 (
            .O(N__32466),
            .I(N__32419));
    Span4Mux_v I__6219 (
            .O(N__32453),
            .I(N__32419));
    Span4Mux_h I__6218 (
            .O(N__32448),
            .I(N__32419));
    Sp12to4 I__6217 (
            .O(N__32443),
            .I(N__32412));
    Sp12to4 I__6216 (
            .O(N__32438),
            .I(N__32412));
    LocalMux I__6215 (
            .O(N__32435),
            .I(N__32412));
    Span4Mux_h I__6214 (
            .O(N__32432),
            .I(N__32409));
    Span4Mux_h I__6213 (
            .O(N__32419),
            .I(N__32406));
    Odrv12 I__6212 (
            .O(N__32412),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__6211 (
            .O(N__32409),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__6210 (
            .O(N__32406),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__6209 (
            .O(N__32399),
            .I(N__32396));
    LocalMux I__6208 (
            .O(N__32396),
            .I(N__32392));
    InMux I__6207 (
            .O(N__32395),
            .I(N__32389));
    Odrv12 I__6206 (
            .O(N__32392),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    LocalMux I__6205 (
            .O(N__32389),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ));
    CascadeMux I__6204 (
            .O(N__32384),
            .I(N__32381));
    InMux I__6203 (
            .O(N__32381),
            .I(N__32378));
    LocalMux I__6202 (
            .O(N__32378),
            .I(N__32374));
    CascadeMux I__6201 (
            .O(N__32377),
            .I(N__32369));
    Span4Mux_h I__6200 (
            .O(N__32374),
            .I(N__32365));
    InMux I__6199 (
            .O(N__32373),
            .I(N__32360));
    InMux I__6198 (
            .O(N__32372),
            .I(N__32360));
    InMux I__6197 (
            .O(N__32369),
            .I(N__32357));
    InMux I__6196 (
            .O(N__32368),
            .I(N__32354));
    Span4Mux_h I__6195 (
            .O(N__32365),
            .I(N__32349));
    LocalMux I__6194 (
            .O(N__32360),
            .I(N__32349));
    LocalMux I__6193 (
            .O(N__32357),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    LocalMux I__6192 (
            .O(N__32354),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__6191 (
            .O(N__32349),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    CascadeMux I__6190 (
            .O(N__32342),
            .I(N__32339));
    InMux I__6189 (
            .O(N__32339),
            .I(N__32336));
    LocalMux I__6188 (
            .O(N__32336),
            .I(N__32332));
    InMux I__6187 (
            .O(N__32335),
            .I(N__32329));
    Span4Mux_v I__6186 (
            .O(N__32332),
            .I(N__32323));
    LocalMux I__6185 (
            .O(N__32329),
            .I(N__32323));
    InMux I__6184 (
            .O(N__32328),
            .I(N__32320));
    Span4Mux_v I__6183 (
            .O(N__32323),
            .I(N__32317));
    LocalMux I__6182 (
            .O(N__32320),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__6181 (
            .O(N__32317),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__6180 (
            .O(N__32312),
            .I(N__32309));
    InMux I__6179 (
            .O(N__32309),
            .I(N__32305));
    InMux I__6178 (
            .O(N__32308),
            .I(N__32302));
    LocalMux I__6177 (
            .O(N__32305),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    LocalMux I__6176 (
            .O(N__32302),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__6175 (
            .O(N__32297),
            .I(N__32287));
    InMux I__6174 (
            .O(N__32296),
            .I(N__32287));
    InMux I__6173 (
            .O(N__32295),
            .I(N__32287));
    CascadeMux I__6172 (
            .O(N__32294),
            .I(N__32283));
    LocalMux I__6171 (
            .O(N__32287),
            .I(N__32280));
    InMux I__6170 (
            .O(N__32286),
            .I(N__32275));
    InMux I__6169 (
            .O(N__32283),
            .I(N__32275));
    Span4Mux_h I__6168 (
            .O(N__32280),
            .I(N__32272));
    LocalMux I__6167 (
            .O(N__32275),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__6166 (
            .O(N__32272),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    InMux I__6165 (
            .O(N__32267),
            .I(N__32263));
    InMux I__6164 (
            .O(N__32266),
            .I(N__32258));
    LocalMux I__6163 (
            .O(N__32263),
            .I(N__32255));
    InMux I__6162 (
            .O(N__32262),
            .I(N__32252));
    CascadeMux I__6161 (
            .O(N__32261),
            .I(N__32249));
    LocalMux I__6160 (
            .O(N__32258),
            .I(N__32242));
    Span4Mux_v I__6159 (
            .O(N__32255),
            .I(N__32242));
    LocalMux I__6158 (
            .O(N__32252),
            .I(N__32242));
    InMux I__6157 (
            .O(N__32249),
            .I(N__32239));
    Span4Mux_v I__6156 (
            .O(N__32242),
            .I(N__32236));
    LocalMux I__6155 (
            .O(N__32239),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__6154 (
            .O(N__32236),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__6153 (
            .O(N__32231),
            .I(N__32225));
    InMux I__6152 (
            .O(N__32230),
            .I(N__32222));
    InMux I__6151 (
            .O(N__32229),
            .I(N__32216));
    InMux I__6150 (
            .O(N__32228),
            .I(N__32216));
    LocalMux I__6149 (
            .O(N__32225),
            .I(N__32213));
    LocalMux I__6148 (
            .O(N__32222),
            .I(N__32210));
    InMux I__6147 (
            .O(N__32221),
            .I(N__32207));
    LocalMux I__6146 (
            .O(N__32216),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv12 I__6145 (
            .O(N__32213),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__6144 (
            .O(N__32210),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__6143 (
            .O(N__32207),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    IoInMux I__6142 (
            .O(N__32198),
            .I(N__32195));
    LocalMux I__6141 (
            .O(N__32195),
            .I(N__32192));
    Span4Mux_s1_v I__6140 (
            .O(N__32192),
            .I(N__32169));
    InMux I__6139 (
            .O(N__32191),
            .I(N__32156));
    InMux I__6138 (
            .O(N__32190),
            .I(N__32156));
    InMux I__6137 (
            .O(N__32189),
            .I(N__32156));
    InMux I__6136 (
            .O(N__32188),
            .I(N__32156));
    InMux I__6135 (
            .O(N__32187),
            .I(N__32147));
    InMux I__6134 (
            .O(N__32186),
            .I(N__32147));
    InMux I__6133 (
            .O(N__32185),
            .I(N__32147));
    InMux I__6132 (
            .O(N__32184),
            .I(N__32147));
    InMux I__6131 (
            .O(N__32183),
            .I(N__32140));
    InMux I__6130 (
            .O(N__32182),
            .I(N__32140));
    InMux I__6129 (
            .O(N__32181),
            .I(N__32140));
    InMux I__6128 (
            .O(N__32180),
            .I(N__32131));
    InMux I__6127 (
            .O(N__32179),
            .I(N__32131));
    InMux I__6126 (
            .O(N__32178),
            .I(N__32131));
    InMux I__6125 (
            .O(N__32177),
            .I(N__32131));
    InMux I__6124 (
            .O(N__32176),
            .I(N__32122));
    InMux I__6123 (
            .O(N__32175),
            .I(N__32122));
    InMux I__6122 (
            .O(N__32174),
            .I(N__32122));
    InMux I__6121 (
            .O(N__32173),
            .I(N__32122));
    InMux I__6120 (
            .O(N__32172),
            .I(N__32119));
    Sp12to4 I__6119 (
            .O(N__32169),
            .I(N__32116));
    InMux I__6118 (
            .O(N__32168),
            .I(N__32100));
    InMux I__6117 (
            .O(N__32167),
            .I(N__32100));
    InMux I__6116 (
            .O(N__32166),
            .I(N__32100));
    InMux I__6115 (
            .O(N__32165),
            .I(N__32100));
    LocalMux I__6114 (
            .O(N__32156),
            .I(N__32097));
    LocalMux I__6113 (
            .O(N__32147),
            .I(N__32086));
    LocalMux I__6112 (
            .O(N__32140),
            .I(N__32086));
    LocalMux I__6111 (
            .O(N__32131),
            .I(N__32086));
    LocalMux I__6110 (
            .O(N__32122),
            .I(N__32086));
    LocalMux I__6109 (
            .O(N__32119),
            .I(N__32086));
    Span12Mux_h I__6108 (
            .O(N__32116),
            .I(N__32083));
    InMux I__6107 (
            .O(N__32115),
            .I(N__32076));
    InMux I__6106 (
            .O(N__32114),
            .I(N__32076));
    InMux I__6105 (
            .O(N__32113),
            .I(N__32076));
    InMux I__6104 (
            .O(N__32112),
            .I(N__32067));
    InMux I__6103 (
            .O(N__32111),
            .I(N__32067));
    InMux I__6102 (
            .O(N__32110),
            .I(N__32067));
    InMux I__6101 (
            .O(N__32109),
            .I(N__32067));
    LocalMux I__6100 (
            .O(N__32100),
            .I(N__32064));
    Span4Mux_v I__6099 (
            .O(N__32097),
            .I(N__32059));
    Span4Mux_v I__6098 (
            .O(N__32086),
            .I(N__32059));
    Span12Mux_v I__6097 (
            .O(N__32083),
            .I(N__32056));
    LocalMux I__6096 (
            .O(N__32076),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    LocalMux I__6095 (
            .O(N__32067),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__6094 (
            .O(N__32064),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__6093 (
            .O(N__32059),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv12 I__6092 (
            .O(N__32056),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__6091 (
            .O(N__32045),
            .I(N__32042));
    LocalMux I__6090 (
            .O(N__32042),
            .I(N__32036));
    InMux I__6089 (
            .O(N__32041),
            .I(N__32033));
    InMux I__6088 (
            .O(N__32040),
            .I(N__32030));
    InMux I__6087 (
            .O(N__32039),
            .I(N__32027));
    Span4Mux_v I__6086 (
            .O(N__32036),
            .I(N__32022));
    LocalMux I__6085 (
            .O(N__32033),
            .I(N__32022));
    LocalMux I__6084 (
            .O(N__32030),
            .I(N__32017));
    LocalMux I__6083 (
            .O(N__32027),
            .I(N__32017));
    Span4Mux_v I__6082 (
            .O(N__32022),
            .I(N__32012));
    Span4Mux_v I__6081 (
            .O(N__32017),
            .I(N__32012));
    Odrv4 I__6080 (
            .O(N__32012),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__6079 (
            .O(N__32009),
            .I(N__32000));
    InMux I__6078 (
            .O(N__32008),
            .I(N__31997));
    InMux I__6077 (
            .O(N__32007),
            .I(N__31960));
    InMux I__6076 (
            .O(N__32006),
            .I(N__31953));
    InMux I__6075 (
            .O(N__32005),
            .I(N__31950));
    InMux I__6074 (
            .O(N__32004),
            .I(N__31947));
    InMux I__6073 (
            .O(N__32003),
            .I(N__31944));
    LocalMux I__6072 (
            .O(N__32000),
            .I(N__31932));
    LocalMux I__6071 (
            .O(N__31997),
            .I(N__31932));
    InMux I__6070 (
            .O(N__31996),
            .I(N__31925));
    InMux I__6069 (
            .O(N__31995),
            .I(N__31925));
    InMux I__6068 (
            .O(N__31994),
            .I(N__31925));
    InMux I__6067 (
            .O(N__31993),
            .I(N__31922));
    InMux I__6066 (
            .O(N__31992),
            .I(N__31913));
    InMux I__6065 (
            .O(N__31991),
            .I(N__31913));
    InMux I__6064 (
            .O(N__31990),
            .I(N__31913));
    InMux I__6063 (
            .O(N__31989),
            .I(N__31913));
    CascadeMux I__6062 (
            .O(N__31988),
            .I(N__31895));
    InMux I__6061 (
            .O(N__31987),
            .I(N__31885));
    InMux I__6060 (
            .O(N__31986),
            .I(N__31885));
    InMux I__6059 (
            .O(N__31985),
            .I(N__31885));
    InMux I__6058 (
            .O(N__31984),
            .I(N__31885));
    InMux I__6057 (
            .O(N__31983),
            .I(N__31882));
    InMux I__6056 (
            .O(N__31982),
            .I(N__31865));
    InMux I__6055 (
            .O(N__31981),
            .I(N__31865));
    InMux I__6054 (
            .O(N__31980),
            .I(N__31865));
    InMux I__6053 (
            .O(N__31979),
            .I(N__31865));
    InMux I__6052 (
            .O(N__31978),
            .I(N__31865));
    InMux I__6051 (
            .O(N__31977),
            .I(N__31865));
    InMux I__6050 (
            .O(N__31976),
            .I(N__31865));
    InMux I__6049 (
            .O(N__31975),
            .I(N__31865));
    InMux I__6048 (
            .O(N__31974),
            .I(N__31854));
    InMux I__6047 (
            .O(N__31973),
            .I(N__31854));
    InMux I__6046 (
            .O(N__31972),
            .I(N__31854));
    InMux I__6045 (
            .O(N__31971),
            .I(N__31854));
    InMux I__6044 (
            .O(N__31970),
            .I(N__31854));
    InMux I__6043 (
            .O(N__31969),
            .I(N__31849));
    InMux I__6042 (
            .O(N__31968),
            .I(N__31849));
    InMux I__6041 (
            .O(N__31967),
            .I(N__31838));
    InMux I__6040 (
            .O(N__31966),
            .I(N__31838));
    InMux I__6039 (
            .O(N__31965),
            .I(N__31838));
    InMux I__6038 (
            .O(N__31964),
            .I(N__31838));
    InMux I__6037 (
            .O(N__31963),
            .I(N__31838));
    LocalMux I__6036 (
            .O(N__31960),
            .I(N__31835));
    InMux I__6035 (
            .O(N__31959),
            .I(N__31830));
    InMux I__6034 (
            .O(N__31958),
            .I(N__31823));
    InMux I__6033 (
            .O(N__31957),
            .I(N__31823));
    InMux I__6032 (
            .O(N__31956),
            .I(N__31823));
    LocalMux I__6031 (
            .O(N__31953),
            .I(N__31816));
    LocalMux I__6030 (
            .O(N__31950),
            .I(N__31816));
    LocalMux I__6029 (
            .O(N__31947),
            .I(N__31816));
    LocalMux I__6028 (
            .O(N__31944),
            .I(N__31809));
    InMux I__6027 (
            .O(N__31943),
            .I(N__31806));
    InMux I__6026 (
            .O(N__31942),
            .I(N__31801));
    InMux I__6025 (
            .O(N__31941),
            .I(N__31801));
    InMux I__6024 (
            .O(N__31940),
            .I(N__31796));
    InMux I__6023 (
            .O(N__31939),
            .I(N__31796));
    InMux I__6022 (
            .O(N__31938),
            .I(N__31793));
    InMux I__6021 (
            .O(N__31937),
            .I(N__31790));
    Span4Mux_h I__6020 (
            .O(N__31932),
            .I(N__31781));
    LocalMux I__6019 (
            .O(N__31925),
            .I(N__31781));
    LocalMux I__6018 (
            .O(N__31922),
            .I(N__31781));
    LocalMux I__6017 (
            .O(N__31913),
            .I(N__31781));
    InMux I__6016 (
            .O(N__31912),
            .I(N__31766));
    InMux I__6015 (
            .O(N__31911),
            .I(N__31761));
    InMux I__6014 (
            .O(N__31910),
            .I(N__31750));
    InMux I__6013 (
            .O(N__31909),
            .I(N__31750));
    InMux I__6012 (
            .O(N__31908),
            .I(N__31750));
    InMux I__6011 (
            .O(N__31907),
            .I(N__31750));
    InMux I__6010 (
            .O(N__31906),
            .I(N__31750));
    InMux I__6009 (
            .O(N__31905),
            .I(N__31743));
    InMux I__6008 (
            .O(N__31904),
            .I(N__31740));
    InMux I__6007 (
            .O(N__31903),
            .I(N__31731));
    InMux I__6006 (
            .O(N__31902),
            .I(N__31731));
    InMux I__6005 (
            .O(N__31901),
            .I(N__31731));
    InMux I__6004 (
            .O(N__31900),
            .I(N__31731));
    InMux I__6003 (
            .O(N__31899),
            .I(N__31722));
    InMux I__6002 (
            .O(N__31898),
            .I(N__31722));
    InMux I__6001 (
            .O(N__31895),
            .I(N__31722));
    InMux I__6000 (
            .O(N__31894),
            .I(N__31722));
    LocalMux I__5999 (
            .O(N__31885),
            .I(N__31719));
    LocalMux I__5998 (
            .O(N__31882),
            .I(N__31706));
    LocalMux I__5997 (
            .O(N__31865),
            .I(N__31706));
    LocalMux I__5996 (
            .O(N__31854),
            .I(N__31706));
    LocalMux I__5995 (
            .O(N__31849),
            .I(N__31706));
    LocalMux I__5994 (
            .O(N__31838),
            .I(N__31706));
    Span4Mux_s3_v I__5993 (
            .O(N__31835),
            .I(N__31706));
    InMux I__5992 (
            .O(N__31834),
            .I(N__31701));
    InMux I__5991 (
            .O(N__31833),
            .I(N__31701));
    LocalMux I__5990 (
            .O(N__31830),
            .I(N__31698));
    LocalMux I__5989 (
            .O(N__31823),
            .I(N__31693));
    Span4Mux_v I__5988 (
            .O(N__31816),
            .I(N__31693));
    InMux I__5987 (
            .O(N__31815),
            .I(N__31684));
    InMux I__5986 (
            .O(N__31814),
            .I(N__31684));
    InMux I__5985 (
            .O(N__31813),
            .I(N__31684));
    InMux I__5984 (
            .O(N__31812),
            .I(N__31684));
    Span4Mux_h I__5983 (
            .O(N__31809),
            .I(N__31679));
    LocalMux I__5982 (
            .O(N__31806),
            .I(N__31679));
    LocalMux I__5981 (
            .O(N__31801),
            .I(N__31674));
    LocalMux I__5980 (
            .O(N__31796),
            .I(N__31674));
    LocalMux I__5979 (
            .O(N__31793),
            .I(N__31671));
    LocalMux I__5978 (
            .O(N__31790),
            .I(N__31668));
    Span4Mux_v I__5977 (
            .O(N__31781),
            .I(N__31665));
    InMux I__5976 (
            .O(N__31780),
            .I(N__31656));
    InMux I__5975 (
            .O(N__31779),
            .I(N__31656));
    InMux I__5974 (
            .O(N__31778),
            .I(N__31656));
    InMux I__5973 (
            .O(N__31777),
            .I(N__31656));
    InMux I__5972 (
            .O(N__31776),
            .I(N__31645));
    InMux I__5971 (
            .O(N__31775),
            .I(N__31645));
    InMux I__5970 (
            .O(N__31774),
            .I(N__31645));
    InMux I__5969 (
            .O(N__31773),
            .I(N__31645));
    InMux I__5968 (
            .O(N__31772),
            .I(N__31645));
    InMux I__5967 (
            .O(N__31771),
            .I(N__31638));
    InMux I__5966 (
            .O(N__31770),
            .I(N__31638));
    InMux I__5965 (
            .O(N__31769),
            .I(N__31638));
    LocalMux I__5964 (
            .O(N__31766),
            .I(N__31635));
    InMux I__5963 (
            .O(N__31765),
            .I(N__31630));
    InMux I__5962 (
            .O(N__31764),
            .I(N__31630));
    LocalMux I__5961 (
            .O(N__31761),
            .I(N__31625));
    LocalMux I__5960 (
            .O(N__31750),
            .I(N__31625));
    InMux I__5959 (
            .O(N__31749),
            .I(N__31616));
    InMux I__5958 (
            .O(N__31748),
            .I(N__31616));
    InMux I__5957 (
            .O(N__31747),
            .I(N__31616));
    InMux I__5956 (
            .O(N__31746),
            .I(N__31616));
    LocalMux I__5955 (
            .O(N__31743),
            .I(N__31603));
    LocalMux I__5954 (
            .O(N__31740),
            .I(N__31603));
    LocalMux I__5953 (
            .O(N__31731),
            .I(N__31603));
    LocalMux I__5952 (
            .O(N__31722),
            .I(N__31603));
    Span4Mux_h I__5951 (
            .O(N__31719),
            .I(N__31603));
    Span4Mux_v I__5950 (
            .O(N__31706),
            .I(N__31603));
    LocalMux I__5949 (
            .O(N__31701),
            .I(N__31584));
    Span4Mux_v I__5948 (
            .O(N__31698),
            .I(N__31584));
    Span4Mux_v I__5947 (
            .O(N__31693),
            .I(N__31584));
    LocalMux I__5946 (
            .O(N__31684),
            .I(N__31584));
    Span4Mux_v I__5945 (
            .O(N__31679),
            .I(N__31584));
    Span4Mux_v I__5944 (
            .O(N__31674),
            .I(N__31584));
    Span4Mux_h I__5943 (
            .O(N__31671),
            .I(N__31584));
    Span4Mux_v I__5942 (
            .O(N__31668),
            .I(N__31584));
    Span4Mux_v I__5941 (
            .O(N__31665),
            .I(N__31584));
    LocalMux I__5940 (
            .O(N__31656),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__5939 (
            .O(N__31645),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__5938 (
            .O(N__31638),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__5937 (
            .O(N__31635),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__5936 (
            .O(N__31630),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__5935 (
            .O(N__31625),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__5934 (
            .O(N__31616),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__5933 (
            .O(N__31603),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__5932 (
            .O(N__31584),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__5931 (
            .O(N__31565),
            .I(N__31562));
    LocalMux I__5930 (
            .O(N__31562),
            .I(N__31557));
    InMux I__5929 (
            .O(N__31561),
            .I(N__31554));
    InMux I__5928 (
            .O(N__31560),
            .I(N__31551));
    Span4Mux_h I__5927 (
            .O(N__31557),
            .I(N__31548));
    LocalMux I__5926 (
            .O(N__31554),
            .I(N__31545));
    LocalMux I__5925 (
            .O(N__31551),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    Odrv4 I__5924 (
            .O(N__31548),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    Odrv12 I__5923 (
            .O(N__31545),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    CascadeMux I__5922 (
            .O(N__31538),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    CascadeMux I__5921 (
            .O(N__31535),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_));
    InMux I__5920 (
            .O(N__31532),
            .I(N__31529));
    LocalMux I__5919 (
            .O(N__31529),
            .I(N__31526));
    Span4Mux_h I__5918 (
            .O(N__31526),
            .I(N__31523));
    Odrv4 I__5917 (
            .O(N__31523),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__5916 (
            .O(N__31520),
            .I(N__31517));
    LocalMux I__5915 (
            .O(N__31517),
            .I(N__31514));
    Odrv12 I__5914 (
            .O(N__31514),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt20 ));
    CascadeMux I__5913 (
            .O(N__31511),
            .I(N__31506));
    InMux I__5912 (
            .O(N__31510),
            .I(N__31503));
    InMux I__5911 (
            .O(N__31509),
            .I(N__31498));
    InMux I__5910 (
            .O(N__31506),
            .I(N__31498));
    LocalMux I__5909 (
            .O(N__31503),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    LocalMux I__5908 (
            .O(N__31498),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    CascadeMux I__5907 (
            .O(N__31493),
            .I(N__31488));
    InMux I__5906 (
            .O(N__31492),
            .I(N__31485));
    InMux I__5905 (
            .O(N__31491),
            .I(N__31480));
    InMux I__5904 (
            .O(N__31488),
            .I(N__31480));
    LocalMux I__5903 (
            .O(N__31485),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    LocalMux I__5902 (
            .O(N__31480),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    CascadeMux I__5901 (
            .O(N__31475),
            .I(N__31472));
    InMux I__5900 (
            .O(N__31472),
            .I(N__31469));
    LocalMux I__5899 (
            .O(N__31469),
            .I(N__31466));
    Odrv4 I__5898 (
            .O(N__31466),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ));
    InMux I__5897 (
            .O(N__31463),
            .I(N__31457));
    InMux I__5896 (
            .O(N__31462),
            .I(N__31457));
    LocalMux I__5895 (
            .O(N__31457),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ));
    InMux I__5894 (
            .O(N__31454),
            .I(N__31450));
    InMux I__5893 (
            .O(N__31453),
            .I(N__31447));
    LocalMux I__5892 (
            .O(N__31450),
            .I(N__31443));
    LocalMux I__5891 (
            .O(N__31447),
            .I(N__31440));
    InMux I__5890 (
            .O(N__31446),
            .I(N__31437));
    Span12Mux_h I__5889 (
            .O(N__31443),
            .I(N__31434));
    Span4Mux_h I__5888 (
            .O(N__31440),
            .I(N__31431));
    LocalMux I__5887 (
            .O(N__31437),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv12 I__5886 (
            .O(N__31434),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv4 I__5885 (
            .O(N__31431),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    InMux I__5884 (
            .O(N__31424),
            .I(N__31421));
    LocalMux I__5883 (
            .O(N__31421),
            .I(N__31417));
    InMux I__5882 (
            .O(N__31420),
            .I(N__31414));
    Span4Mux_v I__5881 (
            .O(N__31417),
            .I(N__31410));
    LocalMux I__5880 (
            .O(N__31414),
            .I(N__31406));
    InMux I__5879 (
            .O(N__31413),
            .I(N__31403));
    Span4Mux_v I__5878 (
            .O(N__31410),
            .I(N__31400));
    InMux I__5877 (
            .O(N__31409),
            .I(N__31397));
    Span4Mux_h I__5876 (
            .O(N__31406),
            .I(N__31392));
    LocalMux I__5875 (
            .O(N__31403),
            .I(N__31392));
    Span4Mux_h I__5874 (
            .O(N__31400),
            .I(N__31387));
    LocalMux I__5873 (
            .O(N__31397),
            .I(N__31387));
    Odrv4 I__5872 (
            .O(N__31392),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv4 I__5871 (
            .O(N__31387),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__5870 (
            .O(N__31382),
            .I(N__31376));
    InMux I__5869 (
            .O(N__31381),
            .I(N__31376));
    LocalMux I__5868 (
            .O(N__31376),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ));
    InMux I__5867 (
            .O(N__31373),
            .I(N__31368));
    InMux I__5866 (
            .O(N__31372),
            .I(N__31363));
    InMux I__5865 (
            .O(N__31371),
            .I(N__31363));
    LocalMux I__5864 (
            .O(N__31368),
            .I(N__31359));
    LocalMux I__5863 (
            .O(N__31363),
            .I(N__31356));
    InMux I__5862 (
            .O(N__31362),
            .I(N__31353));
    Span4Mux_v I__5861 (
            .O(N__31359),
            .I(N__31350));
    Span4Mux_h I__5860 (
            .O(N__31356),
            .I(N__31345));
    LocalMux I__5859 (
            .O(N__31353),
            .I(N__31345));
    Odrv4 I__5858 (
            .O(N__31350),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__5857 (
            .O(N__31345),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__5856 (
            .O(N__31340),
            .I(N__31336));
    InMux I__5855 (
            .O(N__31339),
            .I(N__31333));
    LocalMux I__5854 (
            .O(N__31336),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    LocalMux I__5853 (
            .O(N__31333),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    InMux I__5852 (
            .O(N__31328),
            .I(N__31325));
    LocalMux I__5851 (
            .O(N__31325),
            .I(N__31322));
    Span4Mux_v I__5850 (
            .O(N__31322),
            .I(N__31319));
    Odrv4 I__5849 (
            .O(N__31319),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    CEMux I__5848 (
            .O(N__31316),
            .I(N__31286));
    CEMux I__5847 (
            .O(N__31315),
            .I(N__31286));
    CEMux I__5846 (
            .O(N__31314),
            .I(N__31286));
    CEMux I__5845 (
            .O(N__31313),
            .I(N__31286));
    CEMux I__5844 (
            .O(N__31312),
            .I(N__31286));
    CEMux I__5843 (
            .O(N__31311),
            .I(N__31286));
    CEMux I__5842 (
            .O(N__31310),
            .I(N__31286));
    CEMux I__5841 (
            .O(N__31309),
            .I(N__31286));
    CEMux I__5840 (
            .O(N__31308),
            .I(N__31286));
    CEMux I__5839 (
            .O(N__31307),
            .I(N__31286));
    GlobalMux I__5838 (
            .O(N__31286),
            .I(N__31283));
    gio2CtrlBuf I__5837 (
            .O(N__31283),
            .I(\phase_controller_inst2.stoper_hc.un1_start_g ));
    CascadeMux I__5836 (
            .O(N__31280),
            .I(N__31277));
    InMux I__5835 (
            .O(N__31277),
            .I(N__31271));
    InMux I__5834 (
            .O(N__31276),
            .I(N__31266));
    InMux I__5833 (
            .O(N__31275),
            .I(N__31266));
    InMux I__5832 (
            .O(N__31274),
            .I(N__31263));
    LocalMux I__5831 (
            .O(N__31271),
            .I(N__31258));
    LocalMux I__5830 (
            .O(N__31266),
            .I(N__31258));
    LocalMux I__5829 (
            .O(N__31263),
            .I(\phase_controller_inst2.hc_time_passed ));
    Odrv12 I__5828 (
            .O(N__31258),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__5827 (
            .O(N__31253),
            .I(N__31247));
    InMux I__5826 (
            .O(N__31252),
            .I(N__31247));
    LocalMux I__5825 (
            .O(N__31247),
            .I(N__31244));
    Span4Mux_h I__5824 (
            .O(N__31244),
            .I(N__31241));
    Odrv4 I__5823 (
            .O(N__31241),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__5822 (
            .O(N__31238),
            .I(N__31233));
    InMux I__5821 (
            .O(N__31237),
            .I(N__31228));
    InMux I__5820 (
            .O(N__31236),
            .I(N__31228));
    LocalMux I__5819 (
            .O(N__31233),
            .I(N__31225));
    LocalMux I__5818 (
            .O(N__31228),
            .I(N__31222));
    Span4Mux_h I__5817 (
            .O(N__31225),
            .I(N__31219));
    Span12Mux_h I__5816 (
            .O(N__31222),
            .I(N__31216));
    IoSpan4Mux I__5815 (
            .O(N__31219),
            .I(N__31213));
    Odrv12 I__5814 (
            .O(N__31216),
            .I(il_min_comp2_c));
    Odrv4 I__5813 (
            .O(N__31213),
            .I(il_min_comp2_c));
    InMux I__5812 (
            .O(N__31208),
            .I(N__31205));
    LocalMux I__5811 (
            .O(N__31205),
            .I(N__31200));
    InMux I__5810 (
            .O(N__31204),
            .I(N__31197));
    InMux I__5809 (
            .O(N__31203),
            .I(N__31194));
    Span4Mux_v I__5808 (
            .O(N__31200),
            .I(N__31187));
    LocalMux I__5807 (
            .O(N__31197),
            .I(N__31187));
    LocalMux I__5806 (
            .O(N__31194),
            .I(N__31187));
    Span4Mux_h I__5805 (
            .O(N__31187),
            .I(N__31184));
    Span4Mux_h I__5804 (
            .O(N__31184),
            .I(N__31181));
    Odrv4 I__5803 (
            .O(N__31181),
            .I(il_max_comp2_c));
    InMux I__5802 (
            .O(N__31178),
            .I(N__31175));
    LocalMux I__5801 (
            .O(N__31175),
            .I(N__31170));
    CascadeMux I__5800 (
            .O(N__31174),
            .I(N__31166));
    InMux I__5799 (
            .O(N__31173),
            .I(N__31163));
    Span12Mux_s11_h I__5798 (
            .O(N__31170),
            .I(N__31160));
    InMux I__5797 (
            .O(N__31169),
            .I(N__31157));
    InMux I__5796 (
            .O(N__31166),
            .I(N__31154));
    LocalMux I__5795 (
            .O(N__31163),
            .I(N__31151));
    Span12Mux_v I__5794 (
            .O(N__31160),
            .I(N__31148));
    LocalMux I__5793 (
            .O(N__31157),
            .I(N__31145));
    LocalMux I__5792 (
            .O(N__31154),
            .I(N__31138));
    Span12Mux_s5_v I__5791 (
            .O(N__31151),
            .I(N__31138));
    Span12Mux_v I__5790 (
            .O(N__31148),
            .I(N__31138));
    Odrv4 I__5789 (
            .O(N__31145),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__5788 (
            .O(N__31138),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    InMux I__5787 (
            .O(N__31133),
            .I(N__31129));
    InMux I__5786 (
            .O(N__31132),
            .I(N__31125));
    LocalMux I__5785 (
            .O(N__31129),
            .I(N__31122));
    CascadeMux I__5784 (
            .O(N__31128),
            .I(N__31118));
    LocalMux I__5783 (
            .O(N__31125),
            .I(N__31113));
    Span4Mux_h I__5782 (
            .O(N__31122),
            .I(N__31113));
    InMux I__5781 (
            .O(N__31121),
            .I(N__31110));
    InMux I__5780 (
            .O(N__31118),
            .I(N__31107));
    Span4Mux_v I__5779 (
            .O(N__31113),
            .I(N__31100));
    LocalMux I__5778 (
            .O(N__31110),
            .I(N__31100));
    LocalMux I__5777 (
            .O(N__31107),
            .I(N__31100));
    Odrv4 I__5776 (
            .O(N__31100),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__5775 (
            .O(N__31097),
            .I(N__31093));
    InMux I__5774 (
            .O(N__31096),
            .I(N__31090));
    LocalMux I__5773 (
            .O(N__31093),
            .I(N__31087));
    LocalMux I__5772 (
            .O(N__31090),
            .I(N__31083));
    Span4Mux_h I__5771 (
            .O(N__31087),
            .I(N__31080));
    InMux I__5770 (
            .O(N__31086),
            .I(N__31077));
    Span4Mux_v I__5769 (
            .O(N__31083),
            .I(N__31074));
    Sp12to4 I__5768 (
            .O(N__31080),
            .I(N__31071));
    LocalMux I__5767 (
            .O(N__31077),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    Odrv4 I__5766 (
            .O(N__31074),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    Odrv12 I__5765 (
            .O(N__31071),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    CascadeMux I__5764 (
            .O(N__31064),
            .I(N__31061));
    InMux I__5763 (
            .O(N__31061),
            .I(N__31058));
    LocalMux I__5762 (
            .O(N__31058),
            .I(N__31055));
    Span4Mux_v I__5761 (
            .O(N__31055),
            .I(N__31052));
    Span4Mux_h I__5760 (
            .O(N__31052),
            .I(N__31049));
    Odrv4 I__5759 (
            .O(N__31049),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt28 ));
    InMux I__5758 (
            .O(N__31046),
            .I(N__31043));
    LocalMux I__5757 (
            .O(N__31043),
            .I(N__31040));
    Span4Mux_h I__5756 (
            .O(N__31040),
            .I(N__31036));
    InMux I__5755 (
            .O(N__31039),
            .I(N__31033));
    Odrv4 I__5754 (
            .O(N__31036),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    LocalMux I__5753 (
            .O(N__31033),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    CascadeMux I__5752 (
            .O(N__31028),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_));
    InMux I__5751 (
            .O(N__31025),
            .I(N__31018));
    InMux I__5750 (
            .O(N__31024),
            .I(N__31018));
    InMux I__5749 (
            .O(N__31023),
            .I(N__31015));
    LocalMux I__5748 (
            .O(N__31018),
            .I(N__31012));
    LocalMux I__5747 (
            .O(N__31015),
            .I(N__31006));
    Span4Mux_h I__5746 (
            .O(N__31012),
            .I(N__31006));
    CascadeMux I__5745 (
            .O(N__31011),
            .I(N__31003));
    Span4Mux_v I__5744 (
            .O(N__31006),
            .I(N__31000));
    InMux I__5743 (
            .O(N__31003),
            .I(N__30997));
    Odrv4 I__5742 (
            .O(N__31000),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__5741 (
            .O(N__30997),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__5740 (
            .O(N__30992),
            .I(N__30986));
    InMux I__5739 (
            .O(N__30991),
            .I(N__30986));
    LocalMux I__5738 (
            .O(N__30986),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    InMux I__5737 (
            .O(N__30983),
            .I(N__30976));
    InMux I__5736 (
            .O(N__30982),
            .I(N__30976));
    InMux I__5735 (
            .O(N__30981),
            .I(N__30973));
    LocalMux I__5734 (
            .O(N__30976),
            .I(N__30970));
    LocalMux I__5733 (
            .O(N__30973),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv12 I__5732 (
            .O(N__30970),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    CascadeMux I__5731 (
            .O(N__30965),
            .I(N__30961));
    CascadeMux I__5730 (
            .O(N__30964),
            .I(N__30958));
    InMux I__5729 (
            .O(N__30961),
            .I(N__30952));
    InMux I__5728 (
            .O(N__30958),
            .I(N__30952));
    InMux I__5727 (
            .O(N__30957),
            .I(N__30949));
    LocalMux I__5726 (
            .O(N__30952),
            .I(N__30946));
    LocalMux I__5725 (
            .O(N__30949),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv12 I__5724 (
            .O(N__30946),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__5723 (
            .O(N__30941),
            .I(N__30935));
    InMux I__5722 (
            .O(N__30940),
            .I(N__30935));
    LocalMux I__5721 (
            .O(N__30935),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    InMux I__5720 (
            .O(N__30932),
            .I(N__30929));
    LocalMux I__5719 (
            .O(N__30929),
            .I(N__30926));
    Span4Mux_h I__5718 (
            .O(N__30926),
            .I(N__30923));
    Odrv4 I__5717 (
            .O(N__30923),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ));
    InMux I__5716 (
            .O(N__30920),
            .I(N__30916));
    InMux I__5715 (
            .O(N__30919),
            .I(N__30912));
    LocalMux I__5714 (
            .O(N__30916),
            .I(N__30909));
    InMux I__5713 (
            .O(N__30915),
            .I(N__30906));
    LocalMux I__5712 (
            .O(N__30912),
            .I(N__30903));
    Span4Mux_v I__5711 (
            .O(N__30909),
            .I(N__30900));
    LocalMux I__5710 (
            .O(N__30906),
            .I(N__30895));
    Span4Mux_h I__5709 (
            .O(N__30903),
            .I(N__30895));
    Span4Mux_h I__5708 (
            .O(N__30900),
            .I(N__30890));
    Span4Mux_v I__5707 (
            .O(N__30895),
            .I(N__30890));
    Odrv4 I__5706 (
            .O(N__30890),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__5705 (
            .O(N__30887),
            .I(N__30884));
    LocalMux I__5704 (
            .O(N__30884),
            .I(N__30881));
    Glb2LocalMux I__5703 (
            .O(N__30881),
            .I(N__30878));
    GlobalMux I__5702 (
            .O(N__30878),
            .I(clk_12mhz));
    IoInMux I__5701 (
            .O(N__30875),
            .I(N__30872));
    LocalMux I__5700 (
            .O(N__30872),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__5699 (
            .O(N__30869),
            .I(N__30866));
    LocalMux I__5698 (
            .O(N__30866),
            .I(\phase_controller_inst2.start_timer_tr_RNO_0_0 ));
    InMux I__5697 (
            .O(N__30863),
            .I(N__30858));
    InMux I__5696 (
            .O(N__30862),
            .I(N__30853));
    InMux I__5695 (
            .O(N__30861),
            .I(N__30853));
    LocalMux I__5694 (
            .O(N__30858),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__5693 (
            .O(N__30853),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__5692 (
            .O(N__30848),
            .I(N__30845));
    LocalMux I__5691 (
            .O(N__30845),
            .I(\phase_controller_inst2.start_timer_hc_0_sqmuxa ));
    InMux I__5690 (
            .O(N__30842),
            .I(N__30839));
    LocalMux I__5689 (
            .O(N__30839),
            .I(N__30835));
    InMux I__5688 (
            .O(N__30838),
            .I(N__30832));
    Odrv4 I__5687 (
            .O(N__30835),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    LocalMux I__5686 (
            .O(N__30832),
            .I(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ));
    InMux I__5685 (
            .O(N__30827),
            .I(N__30821));
    InMux I__5684 (
            .O(N__30826),
            .I(N__30821));
    LocalMux I__5683 (
            .O(N__30821),
            .I(N__30818));
    Span4Mux_s3_v I__5682 (
            .O(N__30818),
            .I(N__30815));
    Span4Mux_h I__5681 (
            .O(N__30815),
            .I(N__30812));
    Sp12to4 I__5680 (
            .O(N__30812),
            .I(N__30807));
    InMux I__5679 (
            .O(N__30811),
            .I(N__30804));
    InMux I__5678 (
            .O(N__30810),
            .I(N__30801));
    Span12Mux_v I__5677 (
            .O(N__30807),
            .I(N__30798));
    LocalMux I__5676 (
            .O(N__30804),
            .I(N__30793));
    LocalMux I__5675 (
            .O(N__30801),
            .I(N__30793));
    Span12Mux_v I__5674 (
            .O(N__30798),
            .I(N__30790));
    Span12Mux_h I__5673 (
            .O(N__30793),
            .I(N__30787));
    Span12Mux_h I__5672 (
            .O(N__30790),
            .I(N__30782));
    Span12Mux_v I__5671 (
            .O(N__30787),
            .I(N__30782));
    Odrv12 I__5670 (
            .O(N__30782),
            .I(start_stop_c));
    InMux I__5669 (
            .O(N__30779),
            .I(N__30776));
    LocalMux I__5668 (
            .O(N__30776),
            .I(N__30772));
    InMux I__5667 (
            .O(N__30775),
            .I(N__30769));
    Span4Mux_h I__5666 (
            .O(N__30772),
            .I(N__30762));
    LocalMux I__5665 (
            .O(N__30769),
            .I(N__30762));
    InMux I__5664 (
            .O(N__30768),
            .I(N__30759));
    InMux I__5663 (
            .O(N__30767),
            .I(N__30756));
    Odrv4 I__5662 (
            .O(N__30762),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__5661 (
            .O(N__30759),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__5660 (
            .O(N__30756),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__5659 (
            .O(N__30749),
            .I(N__30746));
    LocalMux I__5658 (
            .O(N__30746),
            .I(N__30741));
    InMux I__5657 (
            .O(N__30745),
            .I(N__30738));
    InMux I__5656 (
            .O(N__30744),
            .I(N__30735));
    Span4Mux_h I__5655 (
            .O(N__30741),
            .I(N__30730));
    LocalMux I__5654 (
            .O(N__30738),
            .I(N__30730));
    LocalMux I__5653 (
            .O(N__30735),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    Odrv4 I__5652 (
            .O(N__30730),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    CascadeMux I__5651 (
            .O(N__30725),
            .I(N__30721));
    InMux I__5650 (
            .O(N__30724),
            .I(N__30716));
    InMux I__5649 (
            .O(N__30721),
            .I(N__30713));
    InMux I__5648 (
            .O(N__30720),
            .I(N__30710));
    InMux I__5647 (
            .O(N__30719),
            .I(N__30707));
    LocalMux I__5646 (
            .O(N__30716),
            .I(N__30702));
    LocalMux I__5645 (
            .O(N__30713),
            .I(N__30702));
    LocalMux I__5644 (
            .O(N__30710),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__5643 (
            .O(N__30707),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__5642 (
            .O(N__30702),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    InMux I__5641 (
            .O(N__30695),
            .I(N__30690));
    InMux I__5640 (
            .O(N__30694),
            .I(N__30685));
    InMux I__5639 (
            .O(N__30693),
            .I(N__30685));
    LocalMux I__5638 (
            .O(N__30690),
            .I(N__30680));
    LocalMux I__5637 (
            .O(N__30685),
            .I(N__30680));
    Odrv4 I__5636 (
            .O(N__30680),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    ClkMux I__5635 (
            .O(N__30677),
            .I(N__30671));
    ClkMux I__5634 (
            .O(N__30676),
            .I(N__30671));
    GlobalMux I__5633 (
            .O(N__30671),
            .I(N__30668));
    gio2CtrlBuf I__5632 (
            .O(N__30668),
            .I(delay_tr_input_c_g));
    InMux I__5631 (
            .O(N__30665),
            .I(N__30660));
    InMux I__5630 (
            .O(N__30664),
            .I(N__30657));
    InMux I__5629 (
            .O(N__30663),
            .I(N__30654));
    LocalMux I__5628 (
            .O(N__30660),
            .I(N__30651));
    LocalMux I__5627 (
            .O(N__30657),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__5626 (
            .O(N__30654),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__5625 (
            .O(N__30651),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__5624 (
            .O(N__30644),
            .I(N__30639));
    InMux I__5623 (
            .O(N__30643),
            .I(N__30636));
    InMux I__5622 (
            .O(N__30642),
            .I(N__30633));
    LocalMux I__5621 (
            .O(N__30639),
            .I(N__30630));
    LocalMux I__5620 (
            .O(N__30636),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__5619 (
            .O(N__30633),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__5618 (
            .O(N__30630),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__5617 (
            .O(N__30623),
            .I(N__30619));
    InMux I__5616 (
            .O(N__30622),
            .I(N__30615));
    LocalMux I__5615 (
            .O(N__30619),
            .I(N__30612));
    InMux I__5614 (
            .O(N__30618),
            .I(N__30609));
    LocalMux I__5613 (
            .O(N__30615),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__5612 (
            .O(N__30612),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__5611 (
            .O(N__30609),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__5610 (
            .O(N__30602),
            .I(N__30599));
    LocalMux I__5609 (
            .O(N__30599),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    CascadeMux I__5608 (
            .O(N__30596),
            .I(N__30592));
    InMux I__5607 (
            .O(N__30595),
            .I(N__30588));
    InMux I__5606 (
            .O(N__30592),
            .I(N__30585));
    InMux I__5605 (
            .O(N__30591),
            .I(N__30582));
    LocalMux I__5604 (
            .O(N__30588),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__5603 (
            .O(N__30585),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    LocalMux I__5602 (
            .O(N__30582),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__5601 (
            .O(N__30575),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__5600 (
            .O(N__30572),
            .I(N__30567));
    InMux I__5599 (
            .O(N__30571),
            .I(N__30564));
    InMux I__5598 (
            .O(N__30570),
            .I(N__30561));
    LocalMux I__5597 (
            .O(N__30567),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__5596 (
            .O(N__30564),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    LocalMux I__5595 (
            .O(N__30561),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__5594 (
            .O(N__30554),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__5593 (
            .O(N__30551),
            .I(N__30541));
    InMux I__5592 (
            .O(N__30550),
            .I(N__30541));
    InMux I__5591 (
            .O(N__30549),
            .I(N__30541));
    InMux I__5590 (
            .O(N__30548),
            .I(N__30538));
    LocalMux I__5589 (
            .O(N__30541),
            .I(N__30535));
    LocalMux I__5588 (
            .O(N__30538),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv12 I__5587 (
            .O(N__30535),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__5586 (
            .O(N__30530),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__5585 (
            .O(N__30527),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__5584 (
            .O(N__30524),
            .I(N__30521));
    LocalMux I__5583 (
            .O(N__30521),
            .I(N__30515));
    InMux I__5582 (
            .O(N__30520),
            .I(N__30510));
    InMux I__5581 (
            .O(N__30519),
            .I(N__30510));
    InMux I__5580 (
            .O(N__30518),
            .I(N__30507));
    Sp12to4 I__5579 (
            .O(N__30515),
            .I(N__30502));
    LocalMux I__5578 (
            .O(N__30510),
            .I(N__30502));
    LocalMux I__5577 (
            .O(N__30507),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    Odrv12 I__5576 (
            .O(N__30502),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__5575 (
            .O(N__30497),
            .I(N__30494));
    LocalMux I__5574 (
            .O(N__30494),
            .I(N__30490));
    InMux I__5573 (
            .O(N__30493),
            .I(N__30487));
    Odrv4 I__5572 (
            .O(N__30490),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    LocalMux I__5571 (
            .O(N__30487),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    InMux I__5570 (
            .O(N__30482),
            .I(N__30479));
    LocalMux I__5569 (
            .O(N__30479),
            .I(N__30476));
    Span4Mux_v I__5568 (
            .O(N__30476),
            .I(N__30473));
    Odrv4 I__5567 (
            .O(N__30473),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__5566 (
            .O(N__30470),
            .I(N__30467));
    LocalMux I__5565 (
            .O(N__30467),
            .I(N__30461));
    InMux I__5564 (
            .O(N__30466),
            .I(N__30458));
    InMux I__5563 (
            .O(N__30465),
            .I(N__30455));
    InMux I__5562 (
            .O(N__30464),
            .I(N__30452));
    Odrv4 I__5561 (
            .O(N__30461),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__5560 (
            .O(N__30458),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__5559 (
            .O(N__30455),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__5558 (
            .O(N__30452),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__5557 (
            .O(N__30443),
            .I(N__30440));
    LocalMux I__5556 (
            .O(N__30440),
            .I(N__30436));
    InMux I__5555 (
            .O(N__30439),
            .I(N__30432));
    Span4Mux_h I__5554 (
            .O(N__30436),
            .I(N__30429));
    InMux I__5553 (
            .O(N__30435),
            .I(N__30426));
    LocalMux I__5552 (
            .O(N__30432),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    Odrv4 I__5551 (
            .O(N__30429),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__5550 (
            .O(N__30426),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    CascadeMux I__5549 (
            .O(N__30419),
            .I(N__30416));
    InMux I__5548 (
            .O(N__30416),
            .I(N__30410));
    InMux I__5547 (
            .O(N__30415),
            .I(N__30410));
    LocalMux I__5546 (
            .O(N__30410),
            .I(N__30406));
    InMux I__5545 (
            .O(N__30409),
            .I(N__30403));
    Span4Mux_h I__5544 (
            .O(N__30406),
            .I(N__30400));
    LocalMux I__5543 (
            .O(N__30403),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__5542 (
            .O(N__30400),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__5541 (
            .O(N__30395),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__5540 (
            .O(N__30392),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__5539 (
            .O(N__30389),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    CascadeMux I__5538 (
            .O(N__30386),
            .I(N__30383));
    InMux I__5537 (
            .O(N__30383),
            .I(N__30377));
    InMux I__5536 (
            .O(N__30382),
            .I(N__30377));
    LocalMux I__5535 (
            .O(N__30377),
            .I(N__30373));
    InMux I__5534 (
            .O(N__30376),
            .I(N__30370));
    Span4Mux_h I__5533 (
            .O(N__30373),
            .I(N__30367));
    LocalMux I__5532 (
            .O(N__30370),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__5531 (
            .O(N__30367),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__5530 (
            .O(N__30362),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__5529 (
            .O(N__30359),
            .I(N__30353));
    InMux I__5528 (
            .O(N__30358),
            .I(N__30353));
    LocalMux I__5527 (
            .O(N__30353),
            .I(N__30349));
    InMux I__5526 (
            .O(N__30352),
            .I(N__30346));
    Span4Mux_h I__5525 (
            .O(N__30349),
            .I(N__30343));
    LocalMux I__5524 (
            .O(N__30346),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__5523 (
            .O(N__30343),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__5522 (
            .O(N__30338),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__5521 (
            .O(N__30335),
            .I(N__30330));
    InMux I__5520 (
            .O(N__30334),
            .I(N__30325));
    InMux I__5519 (
            .O(N__30333),
            .I(N__30325));
    LocalMux I__5518 (
            .O(N__30330),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__5517 (
            .O(N__30325),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__5516 (
            .O(N__30320),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    CascadeMux I__5515 (
            .O(N__30317),
            .I(N__30312));
    InMux I__5514 (
            .O(N__30316),
            .I(N__30309));
    InMux I__5513 (
            .O(N__30315),
            .I(N__30304));
    InMux I__5512 (
            .O(N__30312),
            .I(N__30304));
    LocalMux I__5511 (
            .O(N__30309),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__5510 (
            .O(N__30304),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__5509 (
            .O(N__30299),
            .I(bfn_11_11_0_));
    InMux I__5508 (
            .O(N__30296),
            .I(N__30291));
    InMux I__5507 (
            .O(N__30295),
            .I(N__30288));
    InMux I__5506 (
            .O(N__30294),
            .I(N__30285));
    LocalMux I__5505 (
            .O(N__30291),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__5504 (
            .O(N__30288),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__5503 (
            .O(N__30285),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__5502 (
            .O(N__30278),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    CascadeMux I__5501 (
            .O(N__30275),
            .I(N__30271));
    CascadeMux I__5500 (
            .O(N__30274),
            .I(N__30267));
    InMux I__5499 (
            .O(N__30271),
            .I(N__30264));
    InMux I__5498 (
            .O(N__30270),
            .I(N__30261));
    InMux I__5497 (
            .O(N__30267),
            .I(N__30258));
    LocalMux I__5496 (
            .O(N__30264),
            .I(N__30255));
    LocalMux I__5495 (
            .O(N__30261),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__5494 (
            .O(N__30258),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv4 I__5493 (
            .O(N__30255),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__5492 (
            .O(N__30248),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__5491 (
            .O(N__30245),
            .I(N__30241));
    InMux I__5490 (
            .O(N__30244),
            .I(N__30238));
    LocalMux I__5489 (
            .O(N__30241),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__5488 (
            .O(N__30238),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    InMux I__5487 (
            .O(N__30233),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__5486 (
            .O(N__30230),
            .I(N__30226));
    InMux I__5485 (
            .O(N__30229),
            .I(N__30223));
    LocalMux I__5484 (
            .O(N__30226),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__5483 (
            .O(N__30223),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__5482 (
            .O(N__30218),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__5481 (
            .O(N__30215),
            .I(N__30211));
    InMux I__5480 (
            .O(N__30214),
            .I(N__30208));
    LocalMux I__5479 (
            .O(N__30211),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__5478 (
            .O(N__30208),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    InMux I__5477 (
            .O(N__30203),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__5476 (
            .O(N__30200),
            .I(N__30196));
    InMux I__5475 (
            .O(N__30199),
            .I(N__30193));
    LocalMux I__5474 (
            .O(N__30196),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__5473 (
            .O(N__30193),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__5472 (
            .O(N__30188),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__5471 (
            .O(N__30185),
            .I(N__30181));
    InMux I__5470 (
            .O(N__30184),
            .I(N__30178));
    LocalMux I__5469 (
            .O(N__30181),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__5468 (
            .O(N__30178),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    InMux I__5467 (
            .O(N__30173),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    CascadeMux I__5466 (
            .O(N__30170),
            .I(N__30166));
    InMux I__5465 (
            .O(N__30169),
            .I(N__30161));
    InMux I__5464 (
            .O(N__30166),
            .I(N__30161));
    LocalMux I__5463 (
            .O(N__30161),
            .I(N__30157));
    InMux I__5462 (
            .O(N__30160),
            .I(N__30154));
    Span4Mux_h I__5461 (
            .O(N__30157),
            .I(N__30151));
    LocalMux I__5460 (
            .O(N__30154),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__5459 (
            .O(N__30151),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    InMux I__5458 (
            .O(N__30146),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    CascadeMux I__5457 (
            .O(N__30143),
            .I(N__30140));
    InMux I__5456 (
            .O(N__30140),
            .I(N__30135));
    InMux I__5455 (
            .O(N__30139),
            .I(N__30132));
    InMux I__5454 (
            .O(N__30138),
            .I(N__30129));
    LocalMux I__5453 (
            .O(N__30135),
            .I(N__30124));
    LocalMux I__5452 (
            .O(N__30132),
            .I(N__30124));
    LocalMux I__5451 (
            .O(N__30129),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv12 I__5450 (
            .O(N__30124),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    InMux I__5449 (
            .O(N__30119),
            .I(bfn_11_10_0_));
    InMux I__5448 (
            .O(N__30116),
            .I(N__30110));
    InMux I__5447 (
            .O(N__30115),
            .I(N__30110));
    LocalMux I__5446 (
            .O(N__30110),
            .I(N__30106));
    InMux I__5445 (
            .O(N__30109),
            .I(N__30103));
    Span4Mux_h I__5444 (
            .O(N__30106),
            .I(N__30100));
    LocalMux I__5443 (
            .O(N__30103),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__5442 (
            .O(N__30100),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__5441 (
            .O(N__30095),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    CascadeMux I__5440 (
            .O(N__30092),
            .I(N__30089));
    InMux I__5439 (
            .O(N__30089),
            .I(N__30086));
    LocalMux I__5438 (
            .O(N__30086),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ));
    InMux I__5437 (
            .O(N__30083),
            .I(N__30079));
    InMux I__5436 (
            .O(N__30082),
            .I(N__30076));
    LocalMux I__5435 (
            .O(N__30079),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__5434 (
            .O(N__30076),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__5433 (
            .O(N__30071),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__5432 (
            .O(N__30068),
            .I(N__30064));
    InMux I__5431 (
            .O(N__30067),
            .I(N__30061));
    LocalMux I__5430 (
            .O(N__30064),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__5429 (
            .O(N__30061),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    InMux I__5428 (
            .O(N__30056),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__5427 (
            .O(N__30053),
            .I(N__30049));
    InMux I__5426 (
            .O(N__30052),
            .I(N__30046));
    LocalMux I__5425 (
            .O(N__30049),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__5424 (
            .O(N__30046),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__5423 (
            .O(N__30041),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__5422 (
            .O(N__30038),
            .I(N__30034));
    InMux I__5421 (
            .O(N__30037),
            .I(N__30031));
    LocalMux I__5420 (
            .O(N__30034),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__5419 (
            .O(N__30031),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__5418 (
            .O(N__30026),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__5417 (
            .O(N__30023),
            .I(N__30019));
    InMux I__5416 (
            .O(N__30022),
            .I(N__30016));
    LocalMux I__5415 (
            .O(N__30019),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__5414 (
            .O(N__30016),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__5413 (
            .O(N__30011),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__5412 (
            .O(N__30008),
            .I(N__30004));
    InMux I__5411 (
            .O(N__30007),
            .I(N__30001));
    LocalMux I__5410 (
            .O(N__30004),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__5409 (
            .O(N__30001),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    InMux I__5408 (
            .O(N__29996),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__5407 (
            .O(N__29993),
            .I(N__29989));
    InMux I__5406 (
            .O(N__29992),
            .I(N__29986));
    LocalMux I__5405 (
            .O(N__29989),
            .I(N__29983));
    LocalMux I__5404 (
            .O(N__29986),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__5403 (
            .O(N__29983),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__5402 (
            .O(N__29978),
            .I(bfn_11_9_0_));
    InMux I__5401 (
            .O(N__29975),
            .I(N__29971));
    InMux I__5400 (
            .O(N__29974),
            .I(N__29968));
    LocalMux I__5399 (
            .O(N__29971),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__5398 (
            .O(N__29968),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__5397 (
            .O(N__29963),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    CascadeMux I__5396 (
            .O(N__29960),
            .I(\phase_controller_inst2.stoper_hc.un4_running_df30_cascade_ ));
    InMux I__5395 (
            .O(N__29957),
            .I(N__29954));
    LocalMux I__5394 (
            .O(N__29954),
            .I(N__29951));
    Odrv4 I__5393 (
            .O(N__29951),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ));
    CascadeMux I__5392 (
            .O(N__29948),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__5391 (
            .O(N__29945),
            .I(N__29942));
    InMux I__5390 (
            .O(N__29942),
            .I(N__29939));
    LocalMux I__5389 (
            .O(N__29939),
            .I(N__29936));
    Span4Mux_v I__5388 (
            .O(N__29936),
            .I(N__29932));
    InMux I__5387 (
            .O(N__29935),
            .I(N__29929));
    Odrv4 I__5386 (
            .O(N__29932),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    LocalMux I__5385 (
            .O(N__29929),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    CascadeMux I__5384 (
            .O(N__29924),
            .I(N__29921));
    InMux I__5383 (
            .O(N__29921),
            .I(N__29916));
    InMux I__5382 (
            .O(N__29920),
            .I(N__29911));
    InMux I__5381 (
            .O(N__29919),
            .I(N__29911));
    LocalMux I__5380 (
            .O(N__29916),
            .I(N__29908));
    LocalMux I__5379 (
            .O(N__29911),
            .I(N__29905));
    Span4Mux_v I__5378 (
            .O(N__29908),
            .I(N__29902));
    Span4Mux_v I__5377 (
            .O(N__29905),
            .I(N__29899));
    Odrv4 I__5376 (
            .O(N__29902),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    Odrv4 I__5375 (
            .O(N__29899),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    CascadeMux I__5374 (
            .O(N__29894),
            .I(N__29890));
    CascadeMux I__5373 (
            .O(N__29893),
            .I(N__29886));
    InMux I__5372 (
            .O(N__29890),
            .I(N__29879));
    InMux I__5371 (
            .O(N__29889),
            .I(N__29879));
    InMux I__5370 (
            .O(N__29886),
            .I(N__29879));
    LocalMux I__5369 (
            .O(N__29879),
            .I(N__29876));
    Span4Mux_v I__5368 (
            .O(N__29876),
            .I(N__29873));
    Odrv4 I__5367 (
            .O(N__29873),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    InMux I__5366 (
            .O(N__29870),
            .I(N__29867));
    LocalMux I__5365 (
            .O(N__29867),
            .I(N__29864));
    Odrv4 I__5364 (
            .O(N__29864),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    InMux I__5363 (
            .O(N__29861),
            .I(N__29855));
    InMux I__5362 (
            .O(N__29860),
            .I(N__29855));
    LocalMux I__5361 (
            .O(N__29855),
            .I(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ));
    InMux I__5360 (
            .O(N__29852),
            .I(N__29849));
    LocalMux I__5359 (
            .O(N__29849),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ));
    CascadeMux I__5358 (
            .O(N__29846),
            .I(N__29842));
    CascadeMux I__5357 (
            .O(N__29845),
            .I(N__29839));
    InMux I__5356 (
            .O(N__29842),
            .I(N__29835));
    InMux I__5355 (
            .O(N__29839),
            .I(N__29832));
    InMux I__5354 (
            .O(N__29838),
            .I(N__29829));
    LocalMux I__5353 (
            .O(N__29835),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__5352 (
            .O(N__29832),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__5351 (
            .O(N__29829),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__5350 (
            .O(N__29822),
            .I(N__29818));
    InMux I__5349 (
            .O(N__29821),
            .I(N__29815));
    LocalMux I__5348 (
            .O(N__29818),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__5347 (
            .O(N__29815),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    InMux I__5346 (
            .O(N__29810),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    InMux I__5345 (
            .O(N__29807),
            .I(N__29802));
    InMux I__5344 (
            .O(N__29806),
            .I(N__29799));
    InMux I__5343 (
            .O(N__29805),
            .I(N__29796));
    LocalMux I__5342 (
            .O(N__29802),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__5341 (
            .O(N__29799),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__5340 (
            .O(N__29796),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__5339 (
            .O(N__29789),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__5338 (
            .O(N__29786),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__5337 (
            .O(N__29783),
            .I(bfn_10_25_0_));
    InMux I__5336 (
            .O(N__29780),
            .I(N__29766));
    InMux I__5335 (
            .O(N__29779),
            .I(N__29766));
    InMux I__5334 (
            .O(N__29778),
            .I(N__29757));
    InMux I__5333 (
            .O(N__29777),
            .I(N__29757));
    InMux I__5332 (
            .O(N__29776),
            .I(N__29757));
    InMux I__5331 (
            .O(N__29775),
            .I(N__29757));
    InMux I__5330 (
            .O(N__29774),
            .I(N__29748));
    InMux I__5329 (
            .O(N__29773),
            .I(N__29748));
    InMux I__5328 (
            .O(N__29772),
            .I(N__29748));
    InMux I__5327 (
            .O(N__29771),
            .I(N__29748));
    LocalMux I__5326 (
            .O(N__29766),
            .I(N__29745));
    LocalMux I__5325 (
            .O(N__29757),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__5324 (
            .O(N__29748),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__5323 (
            .O(N__29745),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__5322 (
            .O(N__29738),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__5321 (
            .O(N__29735),
            .I(N__29731));
    InMux I__5320 (
            .O(N__29734),
            .I(N__29727));
    LocalMux I__5319 (
            .O(N__29731),
            .I(N__29724));
    InMux I__5318 (
            .O(N__29730),
            .I(N__29721));
    LocalMux I__5317 (
            .O(N__29727),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    Odrv4 I__5316 (
            .O(N__29724),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    LocalMux I__5315 (
            .O(N__29721),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__5314 (
            .O(N__29714),
            .I(N__29710));
    InMux I__5313 (
            .O(N__29713),
            .I(N__29707));
    LocalMux I__5312 (
            .O(N__29710),
            .I(N__29703));
    LocalMux I__5311 (
            .O(N__29707),
            .I(N__29700));
    InMux I__5310 (
            .O(N__29706),
            .I(N__29697));
    Span4Mux_h I__5309 (
            .O(N__29703),
            .I(N__29693));
    Sp12to4 I__5308 (
            .O(N__29700),
            .I(N__29688));
    LocalMux I__5307 (
            .O(N__29697),
            .I(N__29688));
    CascadeMux I__5306 (
            .O(N__29696),
            .I(N__29685));
    Span4Mux_v I__5305 (
            .O(N__29693),
            .I(N__29682));
    Span12Mux_s5_v I__5304 (
            .O(N__29688),
            .I(N__29679));
    InMux I__5303 (
            .O(N__29685),
            .I(N__29676));
    Odrv4 I__5302 (
            .O(N__29682),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv12 I__5301 (
            .O(N__29679),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__5300 (
            .O(N__29676),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    CascadeMux I__5299 (
            .O(N__29669),
            .I(N__29666));
    InMux I__5298 (
            .O(N__29666),
            .I(N__29663));
    LocalMux I__5297 (
            .O(N__29663),
            .I(N__29660));
    Span4Mux_h I__5296 (
            .O(N__29660),
            .I(N__29657));
    Odrv4 I__5295 (
            .O(N__29657),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    InMux I__5294 (
            .O(N__29654),
            .I(N__29648));
    InMux I__5293 (
            .O(N__29653),
            .I(N__29648));
    LocalMux I__5292 (
            .O(N__29648),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    InMux I__5291 (
            .O(N__29645),
            .I(N__29641));
    InMux I__5290 (
            .O(N__29644),
            .I(N__29638));
    LocalMux I__5289 (
            .O(N__29641),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    LocalMux I__5288 (
            .O(N__29638),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    InMux I__5287 (
            .O(N__29633),
            .I(N__29630));
    LocalMux I__5286 (
            .O(N__29630),
            .I(N__29627));
    Odrv4 I__5285 (
            .O(N__29627),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    InMux I__5284 (
            .O(N__29624),
            .I(N__29621));
    LocalMux I__5283 (
            .O(N__29621),
            .I(N__29616));
    InMux I__5282 (
            .O(N__29620),
            .I(N__29611));
    InMux I__5281 (
            .O(N__29619),
            .I(N__29611));
    Span4Mux_v I__5280 (
            .O(N__29616),
            .I(N__29608));
    LocalMux I__5279 (
            .O(N__29611),
            .I(N__29605));
    Span4Mux_v I__5278 (
            .O(N__29608),
            .I(N__29601));
    Sp12to4 I__5277 (
            .O(N__29605),
            .I(N__29598));
    InMux I__5276 (
            .O(N__29604),
            .I(N__29595));
    Odrv4 I__5275 (
            .O(N__29601),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv12 I__5274 (
            .O(N__29598),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    LocalMux I__5273 (
            .O(N__29595),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__5272 (
            .O(N__29588),
            .I(N__29585));
    LocalMux I__5271 (
            .O(N__29585),
            .I(N__29581));
    InMux I__5270 (
            .O(N__29584),
            .I(N__29578));
    Odrv12 I__5269 (
            .O(N__29581),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    LocalMux I__5268 (
            .O(N__29578),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    InMux I__5267 (
            .O(N__29573),
            .I(N__29570));
    LocalMux I__5266 (
            .O(N__29570),
            .I(N__29567));
    Odrv4 I__5265 (
            .O(N__29567),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__5264 (
            .O(N__29564),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    CascadeMux I__5263 (
            .O(N__29561),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__5262 (
            .O(N__29558),
            .I(N__29553));
    InMux I__5261 (
            .O(N__29557),
            .I(N__29550));
    InMux I__5260 (
            .O(N__29556),
            .I(N__29547));
    LocalMux I__5259 (
            .O(N__29553),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__5258 (
            .O(N__29550),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__5257 (
            .O(N__29547),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__5256 (
            .O(N__29540),
            .I(bfn_10_24_0_));
    InMux I__5255 (
            .O(N__29537),
            .I(N__29532));
    InMux I__5254 (
            .O(N__29536),
            .I(N__29529));
    InMux I__5253 (
            .O(N__29535),
            .I(N__29526));
    LocalMux I__5252 (
            .O(N__29532),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__5251 (
            .O(N__29529),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__5250 (
            .O(N__29526),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__5249 (
            .O(N__29519),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__5248 (
            .O(N__29516),
            .I(N__29511));
    InMux I__5247 (
            .O(N__29515),
            .I(N__29508));
    InMux I__5246 (
            .O(N__29514),
            .I(N__29505));
    LocalMux I__5245 (
            .O(N__29511),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__5244 (
            .O(N__29508),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__5243 (
            .O(N__29505),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__5242 (
            .O(N__29498),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__5241 (
            .O(N__29495),
            .I(N__29490));
    InMux I__5240 (
            .O(N__29494),
            .I(N__29487));
    InMux I__5239 (
            .O(N__29493),
            .I(N__29484));
    LocalMux I__5238 (
            .O(N__29490),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__5237 (
            .O(N__29487),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__5236 (
            .O(N__29484),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__5235 (
            .O(N__29477),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__5234 (
            .O(N__29474),
            .I(N__29469));
    InMux I__5233 (
            .O(N__29473),
            .I(N__29466));
    InMux I__5232 (
            .O(N__29472),
            .I(N__29463));
    LocalMux I__5231 (
            .O(N__29469),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__5230 (
            .O(N__29466),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__5229 (
            .O(N__29463),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__5228 (
            .O(N__29456),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__5227 (
            .O(N__29453),
            .I(N__29448));
    InMux I__5226 (
            .O(N__29452),
            .I(N__29445));
    InMux I__5225 (
            .O(N__29451),
            .I(N__29442));
    LocalMux I__5224 (
            .O(N__29448),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__5223 (
            .O(N__29445),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__5222 (
            .O(N__29442),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__5221 (
            .O(N__29435),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__5220 (
            .O(N__29432),
            .I(N__29429));
    LocalMux I__5219 (
            .O(N__29429),
            .I(N__29425));
    InMux I__5218 (
            .O(N__29428),
            .I(N__29421));
    Span4Mux_h I__5217 (
            .O(N__29425),
            .I(N__29418));
    InMux I__5216 (
            .O(N__29424),
            .I(N__29415));
    LocalMux I__5215 (
            .O(N__29421),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    Odrv4 I__5214 (
            .O(N__29418),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    LocalMux I__5213 (
            .O(N__29415),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    InMux I__5212 (
            .O(N__29408),
            .I(N__29404));
    InMux I__5211 (
            .O(N__29407),
            .I(N__29401));
    LocalMux I__5210 (
            .O(N__29404),
            .I(N__29397));
    LocalMux I__5209 (
            .O(N__29401),
            .I(N__29393));
    InMux I__5208 (
            .O(N__29400),
            .I(N__29390));
    Span4Mux_v I__5207 (
            .O(N__29397),
            .I(N__29387));
    InMux I__5206 (
            .O(N__29396),
            .I(N__29384));
    Span4Mux_v I__5205 (
            .O(N__29393),
            .I(N__29379));
    LocalMux I__5204 (
            .O(N__29390),
            .I(N__29379));
    Odrv4 I__5203 (
            .O(N__29387),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    LocalMux I__5202 (
            .O(N__29384),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__5201 (
            .O(N__29379),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    CascadeMux I__5200 (
            .O(N__29372),
            .I(N__29369));
    InMux I__5199 (
            .O(N__29369),
            .I(N__29366));
    LocalMux I__5198 (
            .O(N__29366),
            .I(N__29363));
    Span12Mux_v I__5197 (
            .O(N__29363),
            .I(N__29360));
    Odrv12 I__5196 (
            .O(N__29360),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    CEMux I__5195 (
            .O(N__29357),
            .I(N__29353));
    CEMux I__5194 (
            .O(N__29356),
            .I(N__29350));
    LocalMux I__5193 (
            .O(N__29353),
            .I(N__29345));
    LocalMux I__5192 (
            .O(N__29350),
            .I(N__29342));
    CEMux I__5191 (
            .O(N__29349),
            .I(N__29339));
    CEMux I__5190 (
            .O(N__29348),
            .I(N__29336));
    Span4Mux_v I__5189 (
            .O(N__29345),
            .I(N__29331));
    Span4Mux_v I__5188 (
            .O(N__29342),
            .I(N__29331));
    LocalMux I__5187 (
            .O(N__29339),
            .I(N__29326));
    LocalMux I__5186 (
            .O(N__29336),
            .I(N__29326));
    Span4Mux_h I__5185 (
            .O(N__29331),
            .I(N__29321));
    Span4Mux_v I__5184 (
            .O(N__29326),
            .I(N__29321));
    Odrv4 I__5183 (
            .O(N__29321),
            .I(\delay_measurement_inst.delay_hc_timer.N_203_i ));
    InMux I__5182 (
            .O(N__29318),
            .I(N__29315));
    LocalMux I__5181 (
            .O(N__29315),
            .I(N__29312));
    Span4Mux_h I__5180 (
            .O(N__29312),
            .I(N__29309));
    Sp12to4 I__5179 (
            .O(N__29309),
            .I(N__29306));
    Span12Mux_v I__5178 (
            .O(N__29306),
            .I(N__29303));
    Odrv12 I__5177 (
            .O(N__29303),
            .I(il_max_comp1_D1));
    InMux I__5176 (
            .O(N__29300),
            .I(N__29296));
    InMux I__5175 (
            .O(N__29299),
            .I(N__29293));
    LocalMux I__5174 (
            .O(N__29296),
            .I(N__29290));
    LocalMux I__5173 (
            .O(N__29293),
            .I(N__29287));
    Span4Mux_h I__5172 (
            .O(N__29290),
            .I(N__29282));
    Span4Mux_v I__5171 (
            .O(N__29287),
            .I(N__29282));
    Odrv4 I__5170 (
            .O(N__29282),
            .I(\current_shift_inst.control_input_axb_0 ));
    InMux I__5169 (
            .O(N__29279),
            .I(N__29271));
    InMux I__5168 (
            .O(N__29278),
            .I(N__29271));
    InMux I__5167 (
            .O(N__29277),
            .I(N__29268));
    InMux I__5166 (
            .O(N__29276),
            .I(N__29265));
    LocalMux I__5165 (
            .O(N__29271),
            .I(N__29262));
    LocalMux I__5164 (
            .O(N__29268),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__5163 (
            .O(N__29265),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__5162 (
            .O(N__29262),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__5161 (
            .O(N__29255),
            .I(N__29239));
    InMux I__5160 (
            .O(N__29254),
            .I(N__29239));
    InMux I__5159 (
            .O(N__29253),
            .I(N__29239));
    InMux I__5158 (
            .O(N__29252),
            .I(N__29239));
    InMux I__5157 (
            .O(N__29251),
            .I(N__29208));
    InMux I__5156 (
            .O(N__29250),
            .I(N__29208));
    InMux I__5155 (
            .O(N__29249),
            .I(N__29208));
    InMux I__5154 (
            .O(N__29248),
            .I(N__29208));
    LocalMux I__5153 (
            .O(N__29239),
            .I(N__29205));
    InMux I__5152 (
            .O(N__29238),
            .I(N__29196));
    InMux I__5151 (
            .O(N__29237),
            .I(N__29196));
    InMux I__5150 (
            .O(N__29236),
            .I(N__29196));
    InMux I__5149 (
            .O(N__29235),
            .I(N__29196));
    InMux I__5148 (
            .O(N__29234),
            .I(N__29191));
    InMux I__5147 (
            .O(N__29233),
            .I(N__29191));
    InMux I__5146 (
            .O(N__29232),
            .I(N__29182));
    InMux I__5145 (
            .O(N__29231),
            .I(N__29182));
    InMux I__5144 (
            .O(N__29230),
            .I(N__29182));
    InMux I__5143 (
            .O(N__29229),
            .I(N__29182));
    InMux I__5142 (
            .O(N__29228),
            .I(N__29173));
    InMux I__5141 (
            .O(N__29227),
            .I(N__29173));
    InMux I__5140 (
            .O(N__29226),
            .I(N__29173));
    InMux I__5139 (
            .O(N__29225),
            .I(N__29173));
    InMux I__5138 (
            .O(N__29224),
            .I(N__29164));
    InMux I__5137 (
            .O(N__29223),
            .I(N__29164));
    InMux I__5136 (
            .O(N__29222),
            .I(N__29164));
    InMux I__5135 (
            .O(N__29221),
            .I(N__29164));
    InMux I__5134 (
            .O(N__29220),
            .I(N__29155));
    InMux I__5133 (
            .O(N__29219),
            .I(N__29155));
    InMux I__5132 (
            .O(N__29218),
            .I(N__29155));
    InMux I__5131 (
            .O(N__29217),
            .I(N__29155));
    LocalMux I__5130 (
            .O(N__29208),
            .I(N__29150));
    Span4Mux_v I__5129 (
            .O(N__29205),
            .I(N__29150));
    LocalMux I__5128 (
            .O(N__29196),
            .I(N__29147));
    LocalMux I__5127 (
            .O(N__29191),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__5126 (
            .O(N__29182),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__5125 (
            .O(N__29173),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__5124 (
            .O(N__29164),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    LocalMux I__5123 (
            .O(N__29155),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__5122 (
            .O(N__29150),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__5121 (
            .O(N__29147),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__5120 (
            .O(N__29132),
            .I(N__29129));
    LocalMux I__5119 (
            .O(N__29129),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__5118 (
            .O(N__29126),
            .I(N__29123));
    LocalMux I__5117 (
            .O(N__29123),
            .I(N__29119));
    CascadeMux I__5116 (
            .O(N__29122),
            .I(N__29115));
    Span4Mux_v I__5115 (
            .O(N__29119),
            .I(N__29112));
    InMux I__5114 (
            .O(N__29118),
            .I(N__29109));
    InMux I__5113 (
            .O(N__29115),
            .I(N__29106));
    Odrv4 I__5112 (
            .O(N__29112),
            .I(\current_shift_inst.N_1304_i ));
    LocalMux I__5111 (
            .O(N__29109),
            .I(\current_shift_inst.N_1304_i ));
    LocalMux I__5110 (
            .O(N__29106),
            .I(\current_shift_inst.N_1304_i ));
    CascadeMux I__5109 (
            .O(N__29099),
            .I(N__29096));
    InMux I__5108 (
            .O(N__29096),
            .I(N__29091));
    InMux I__5107 (
            .O(N__29095),
            .I(N__29088));
    InMux I__5106 (
            .O(N__29094),
            .I(N__29085));
    LocalMux I__5105 (
            .O(N__29091),
            .I(N__29080));
    LocalMux I__5104 (
            .O(N__29088),
            .I(N__29080));
    LocalMux I__5103 (
            .O(N__29085),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv4 I__5102 (
            .O(N__29080),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__5101 (
            .O(N__29075),
            .I(N__29071));
    InMux I__5100 (
            .O(N__29074),
            .I(N__29068));
    LocalMux I__5099 (
            .O(N__29071),
            .I(N__29065));
    LocalMux I__5098 (
            .O(N__29068),
            .I(N__29062));
    Span4Mux_h I__5097 (
            .O(N__29065),
            .I(N__29057));
    Span4Mux_v I__5096 (
            .O(N__29062),
            .I(N__29057));
    Span4Mux_v I__5095 (
            .O(N__29057),
            .I(N__29052));
    InMux I__5094 (
            .O(N__29056),
            .I(N__29049));
    InMux I__5093 (
            .O(N__29055),
            .I(N__29046));
    Odrv4 I__5092 (
            .O(N__29052),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__5091 (
            .O(N__29049),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__5090 (
            .O(N__29046),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__5089 (
            .O(N__29039),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__5088 (
            .O(N__29036),
            .I(N__29033));
    InMux I__5087 (
            .O(N__29033),
            .I(N__29029));
    InMux I__5086 (
            .O(N__29032),
            .I(N__29026));
    LocalMux I__5085 (
            .O(N__29029),
            .I(N__29020));
    LocalMux I__5084 (
            .O(N__29026),
            .I(N__29020));
    InMux I__5083 (
            .O(N__29025),
            .I(N__29017));
    Span4Mux_h I__5082 (
            .O(N__29020),
            .I(N__29014));
    LocalMux I__5081 (
            .O(N__29017),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__5080 (
            .O(N__29014),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__5079 (
            .O(N__29009),
            .I(N__29004));
    InMux I__5078 (
            .O(N__29008),
            .I(N__29001));
    InMux I__5077 (
            .O(N__29007),
            .I(N__28998));
    LocalMux I__5076 (
            .O(N__29004),
            .I(N__28995));
    LocalMux I__5075 (
            .O(N__29001),
            .I(N__28992));
    LocalMux I__5074 (
            .O(N__28998),
            .I(N__28989));
    Span4Mux_h I__5073 (
            .O(N__28995),
            .I(N__28984));
    Span4Mux_h I__5072 (
            .O(N__28992),
            .I(N__28984));
    Span12Mux_s10_h I__5071 (
            .O(N__28989),
            .I(N__28978));
    Sp12to4 I__5070 (
            .O(N__28984),
            .I(N__28978));
    InMux I__5069 (
            .O(N__28983),
            .I(N__28975));
    Odrv12 I__5068 (
            .O(N__28978),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    LocalMux I__5067 (
            .O(N__28975),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__5066 (
            .O(N__28970),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__5065 (
            .O(N__28967),
            .I(N__28964));
    InMux I__5064 (
            .O(N__28964),
            .I(N__28960));
    InMux I__5063 (
            .O(N__28963),
            .I(N__28957));
    LocalMux I__5062 (
            .O(N__28960),
            .I(N__28951));
    LocalMux I__5061 (
            .O(N__28957),
            .I(N__28951));
    InMux I__5060 (
            .O(N__28956),
            .I(N__28948));
    Span4Mux_h I__5059 (
            .O(N__28951),
            .I(N__28945));
    LocalMux I__5058 (
            .O(N__28948),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__5057 (
            .O(N__28945),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__5056 (
            .O(N__28940),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__5055 (
            .O(N__28937),
            .I(N__28934));
    InMux I__5054 (
            .O(N__28934),
            .I(N__28930));
    InMux I__5053 (
            .O(N__28933),
            .I(N__28927));
    LocalMux I__5052 (
            .O(N__28930),
            .I(N__28923));
    LocalMux I__5051 (
            .O(N__28927),
            .I(N__28920));
    InMux I__5050 (
            .O(N__28926),
            .I(N__28917));
    Span4Mux_h I__5049 (
            .O(N__28923),
            .I(N__28914));
    Span4Mux_h I__5048 (
            .O(N__28920),
            .I(N__28911));
    LocalMux I__5047 (
            .O(N__28917),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__5046 (
            .O(N__28914),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__5045 (
            .O(N__28911),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__5044 (
            .O(N__28904),
            .I(N__28896));
    InMux I__5043 (
            .O(N__28903),
            .I(N__28896));
    InMux I__5042 (
            .O(N__28902),
            .I(N__28893));
    InMux I__5041 (
            .O(N__28901),
            .I(N__28890));
    LocalMux I__5040 (
            .O(N__28896),
            .I(N__28885));
    LocalMux I__5039 (
            .O(N__28893),
            .I(N__28885));
    LocalMux I__5038 (
            .O(N__28890),
            .I(N__28882));
    Span4Mux_h I__5037 (
            .O(N__28885),
            .I(N__28879));
    Odrv12 I__5036 (
            .O(N__28882),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__5035 (
            .O(N__28879),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__5034 (
            .O(N__28874),
            .I(bfn_10_15_0_));
    InMux I__5033 (
            .O(N__28871),
            .I(N__28867));
    InMux I__5032 (
            .O(N__28870),
            .I(N__28864));
    LocalMux I__5031 (
            .O(N__28867),
            .I(N__28860));
    LocalMux I__5030 (
            .O(N__28864),
            .I(N__28857));
    InMux I__5029 (
            .O(N__28863),
            .I(N__28854));
    Span4Mux_h I__5028 (
            .O(N__28860),
            .I(N__28851));
    Odrv4 I__5027 (
            .O(N__28857),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__5026 (
            .O(N__28854),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__5025 (
            .O(N__28851),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__5024 (
            .O(N__28844),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__5023 (
            .O(N__28841),
            .I(N__28834));
    InMux I__5022 (
            .O(N__28840),
            .I(N__28834));
    InMux I__5021 (
            .O(N__28839),
            .I(N__28831));
    LocalMux I__5020 (
            .O(N__28834),
            .I(N__28828));
    LocalMux I__5019 (
            .O(N__28831),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv4 I__5018 (
            .O(N__28828),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    CascadeMux I__5017 (
            .O(N__28823),
            .I(N__28820));
    InMux I__5016 (
            .O(N__28820),
            .I(N__28816));
    InMux I__5015 (
            .O(N__28819),
            .I(N__28813));
    LocalMux I__5014 (
            .O(N__28816),
            .I(N__28810));
    LocalMux I__5013 (
            .O(N__28813),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv4 I__5012 (
            .O(N__28810),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__5011 (
            .O(N__28805),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__5010 (
            .O(N__28802),
            .I(N__28799));
    LocalMux I__5009 (
            .O(N__28799),
            .I(N__28795));
    InMux I__5008 (
            .O(N__28798),
            .I(N__28792));
    Span4Mux_v I__5007 (
            .O(N__28795),
            .I(N__28789));
    LocalMux I__5006 (
            .O(N__28792),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv4 I__5005 (
            .O(N__28789),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__5004 (
            .O(N__28784),
            .I(N__28779));
    CascadeMux I__5003 (
            .O(N__28783),
            .I(N__28776));
    InMux I__5002 (
            .O(N__28782),
            .I(N__28773));
    InMux I__5001 (
            .O(N__28779),
            .I(N__28768));
    InMux I__5000 (
            .O(N__28776),
            .I(N__28768));
    LocalMux I__4999 (
            .O(N__28773),
            .I(N__28763));
    LocalMux I__4998 (
            .O(N__28768),
            .I(N__28763));
    Odrv4 I__4997 (
            .O(N__28763),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__4996 (
            .O(N__28760),
            .I(N__28755));
    InMux I__4995 (
            .O(N__28759),
            .I(N__28752));
    CascadeMux I__4994 (
            .O(N__28758),
            .I(N__28749));
    LocalMux I__4993 (
            .O(N__28755),
            .I(N__28746));
    LocalMux I__4992 (
            .O(N__28752),
            .I(N__28743));
    InMux I__4991 (
            .O(N__28749),
            .I(N__28740));
    Span4Mux_h I__4990 (
            .O(N__28746),
            .I(N__28732));
    Span4Mux_h I__4989 (
            .O(N__28743),
            .I(N__28732));
    LocalMux I__4988 (
            .O(N__28740),
            .I(N__28732));
    InMux I__4987 (
            .O(N__28739),
            .I(N__28729));
    Odrv4 I__4986 (
            .O(N__28732),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    LocalMux I__4985 (
            .O(N__28729),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__4984 (
            .O(N__28724),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__4983 (
            .O(N__28721),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__4982 (
            .O(N__28718),
            .I(N__28714));
    InMux I__4981 (
            .O(N__28717),
            .I(N__28711));
    LocalMux I__4980 (
            .O(N__28714),
            .I(N__28706));
    LocalMux I__4979 (
            .O(N__28711),
            .I(N__28703));
    InMux I__4978 (
            .O(N__28710),
            .I(N__28698));
    InMux I__4977 (
            .O(N__28709),
            .I(N__28698));
    Span4Mux_h I__4976 (
            .O(N__28706),
            .I(N__28695));
    Span4Mux_v I__4975 (
            .O(N__28703),
            .I(N__28690));
    LocalMux I__4974 (
            .O(N__28698),
            .I(N__28690));
    Odrv4 I__4973 (
            .O(N__28695),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__4972 (
            .O(N__28690),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    CEMux I__4971 (
            .O(N__28685),
            .I(N__28680));
    CEMux I__4970 (
            .O(N__28684),
            .I(N__28677));
    CEMux I__4969 (
            .O(N__28683),
            .I(N__28672));
    LocalMux I__4968 (
            .O(N__28680),
            .I(N__28668));
    LocalMux I__4967 (
            .O(N__28677),
            .I(N__28665));
    CEMux I__4966 (
            .O(N__28676),
            .I(N__28662));
    CEMux I__4965 (
            .O(N__28675),
            .I(N__28659));
    LocalMux I__4964 (
            .O(N__28672),
            .I(N__28656));
    CEMux I__4963 (
            .O(N__28671),
            .I(N__28653));
    Span4Mux_v I__4962 (
            .O(N__28668),
            .I(N__28650));
    Span4Mux_h I__4961 (
            .O(N__28665),
            .I(N__28645));
    LocalMux I__4960 (
            .O(N__28662),
            .I(N__28645));
    LocalMux I__4959 (
            .O(N__28659),
            .I(N__28638));
    Span4Mux_v I__4958 (
            .O(N__28656),
            .I(N__28638));
    LocalMux I__4957 (
            .O(N__28653),
            .I(N__28638));
    Span4Mux_h I__4956 (
            .O(N__28650),
            .I(N__28633));
    Span4Mux_v I__4955 (
            .O(N__28645),
            .I(N__28633));
    Span4Mux_h I__4954 (
            .O(N__28638),
            .I(N__28630));
    Odrv4 I__4953 (
            .O(N__28633),
            .I(\delay_measurement_inst.delay_hc_timer.N_202_i ));
    Odrv4 I__4952 (
            .O(N__28630),
            .I(\delay_measurement_inst.delay_hc_timer.N_202_i ));
    CascadeMux I__4951 (
            .O(N__28625),
            .I(N__28621));
    CascadeMux I__4950 (
            .O(N__28624),
            .I(N__28618));
    InMux I__4949 (
            .O(N__28621),
            .I(N__28612));
    InMux I__4948 (
            .O(N__28618),
            .I(N__28612));
    InMux I__4947 (
            .O(N__28617),
            .I(N__28609));
    LocalMux I__4946 (
            .O(N__28612),
            .I(N__28606));
    LocalMux I__4945 (
            .O(N__28609),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__4944 (
            .O(N__28606),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__4943 (
            .O(N__28601),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__4942 (
            .O(N__28598),
            .I(N__28595));
    InMux I__4941 (
            .O(N__28595),
            .I(N__28591));
    InMux I__4940 (
            .O(N__28594),
            .I(N__28588));
    LocalMux I__4939 (
            .O(N__28591),
            .I(N__28582));
    LocalMux I__4938 (
            .O(N__28588),
            .I(N__28582));
    InMux I__4937 (
            .O(N__28587),
            .I(N__28579));
    Span4Mux_h I__4936 (
            .O(N__28582),
            .I(N__28576));
    LocalMux I__4935 (
            .O(N__28579),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__4934 (
            .O(N__28576),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__4933 (
            .O(N__28571),
            .I(N__28566));
    InMux I__4932 (
            .O(N__28570),
            .I(N__28563));
    InMux I__4931 (
            .O(N__28569),
            .I(N__28560));
    LocalMux I__4930 (
            .O(N__28566),
            .I(N__28557));
    LocalMux I__4929 (
            .O(N__28563),
            .I(N__28552));
    LocalMux I__4928 (
            .O(N__28560),
            .I(N__28552));
    Span4Mux_v I__4927 (
            .O(N__28557),
            .I(N__28547));
    Span4Mux_v I__4926 (
            .O(N__28552),
            .I(N__28547));
    Span4Mux_v I__4925 (
            .O(N__28547),
            .I(N__28543));
    InMux I__4924 (
            .O(N__28546),
            .I(N__28540));
    Odrv4 I__4923 (
            .O(N__28543),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__4922 (
            .O(N__28540),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__4921 (
            .O(N__28535),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__4920 (
            .O(N__28532),
            .I(N__28529));
    InMux I__4919 (
            .O(N__28529),
            .I(N__28525));
    InMux I__4918 (
            .O(N__28528),
            .I(N__28522));
    LocalMux I__4917 (
            .O(N__28525),
            .I(N__28516));
    LocalMux I__4916 (
            .O(N__28522),
            .I(N__28516));
    InMux I__4915 (
            .O(N__28521),
            .I(N__28513));
    Span4Mux_h I__4914 (
            .O(N__28516),
            .I(N__28510));
    LocalMux I__4913 (
            .O(N__28513),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__4912 (
            .O(N__28510),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__4911 (
            .O(N__28505),
            .I(N__28500));
    InMux I__4910 (
            .O(N__28504),
            .I(N__28495));
    InMux I__4909 (
            .O(N__28503),
            .I(N__28495));
    LocalMux I__4908 (
            .O(N__28500),
            .I(N__28492));
    LocalMux I__4907 (
            .O(N__28495),
            .I(N__28489));
    Span4Mux_h I__4906 (
            .O(N__28492),
            .I(N__28484));
    Span4Mux_h I__4905 (
            .O(N__28489),
            .I(N__28484));
    Span4Mux_v I__4904 (
            .O(N__28484),
            .I(N__28480));
    InMux I__4903 (
            .O(N__28483),
            .I(N__28477));
    Odrv4 I__4902 (
            .O(N__28480),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__4901 (
            .O(N__28477),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__4900 (
            .O(N__28472),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__4899 (
            .O(N__28469),
            .I(N__28466));
    InMux I__4898 (
            .O(N__28466),
            .I(N__28462));
    InMux I__4897 (
            .O(N__28465),
            .I(N__28459));
    LocalMux I__4896 (
            .O(N__28462),
            .I(N__28455));
    LocalMux I__4895 (
            .O(N__28459),
            .I(N__28452));
    InMux I__4894 (
            .O(N__28458),
            .I(N__28449));
    Span4Mux_h I__4893 (
            .O(N__28455),
            .I(N__28446));
    Span4Mux_h I__4892 (
            .O(N__28452),
            .I(N__28443));
    LocalMux I__4891 (
            .O(N__28449),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__4890 (
            .O(N__28446),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__4889 (
            .O(N__28443),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__4888 (
            .O(N__28436),
            .I(N__28430));
    InMux I__4887 (
            .O(N__28435),
            .I(N__28427));
    CascadeMux I__4886 (
            .O(N__28434),
            .I(N__28424));
    InMux I__4885 (
            .O(N__28433),
            .I(N__28421));
    LocalMux I__4884 (
            .O(N__28430),
            .I(N__28418));
    LocalMux I__4883 (
            .O(N__28427),
            .I(N__28415));
    InMux I__4882 (
            .O(N__28424),
            .I(N__28412));
    LocalMux I__4881 (
            .O(N__28421),
            .I(N__28409));
    Span4Mux_v I__4880 (
            .O(N__28418),
            .I(N__28404));
    Span4Mux_h I__4879 (
            .O(N__28415),
            .I(N__28404));
    LocalMux I__4878 (
            .O(N__28412),
            .I(N__28401));
    Span4Mux_v I__4877 (
            .O(N__28409),
            .I(N__28396));
    Span4Mux_v I__4876 (
            .O(N__28404),
            .I(N__28396));
    Span4Mux_h I__4875 (
            .O(N__28401),
            .I(N__28393));
    Odrv4 I__4874 (
            .O(N__28396),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    Odrv4 I__4873 (
            .O(N__28393),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__4872 (
            .O(N__28388),
            .I(bfn_10_14_0_));
    InMux I__4871 (
            .O(N__28385),
            .I(N__28381));
    InMux I__4870 (
            .O(N__28384),
            .I(N__28378));
    LocalMux I__4869 (
            .O(N__28381),
            .I(N__28374));
    LocalMux I__4868 (
            .O(N__28378),
            .I(N__28371));
    InMux I__4867 (
            .O(N__28377),
            .I(N__28368));
    Span4Mux_h I__4866 (
            .O(N__28374),
            .I(N__28365));
    Span4Mux_h I__4865 (
            .O(N__28371),
            .I(N__28362));
    LocalMux I__4864 (
            .O(N__28368),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__4863 (
            .O(N__28365),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__4862 (
            .O(N__28362),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__4861 (
            .O(N__28355),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__4860 (
            .O(N__28352),
            .I(N__28345));
    InMux I__4859 (
            .O(N__28351),
            .I(N__28345));
    InMux I__4858 (
            .O(N__28350),
            .I(N__28342));
    LocalMux I__4857 (
            .O(N__28345),
            .I(N__28339));
    LocalMux I__4856 (
            .O(N__28342),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__4855 (
            .O(N__28339),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__4854 (
            .O(N__28334),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__4853 (
            .O(N__28331),
            .I(N__28327));
    CascadeMux I__4852 (
            .O(N__28330),
            .I(N__28324));
    InMux I__4851 (
            .O(N__28327),
            .I(N__28318));
    InMux I__4850 (
            .O(N__28324),
            .I(N__28318));
    InMux I__4849 (
            .O(N__28323),
            .I(N__28315));
    LocalMux I__4848 (
            .O(N__28318),
            .I(N__28312));
    LocalMux I__4847 (
            .O(N__28315),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv4 I__4846 (
            .O(N__28312),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__4845 (
            .O(N__28307),
            .I(N__28302));
    InMux I__4844 (
            .O(N__28306),
            .I(N__28297));
    InMux I__4843 (
            .O(N__28305),
            .I(N__28297));
    LocalMux I__4842 (
            .O(N__28302),
            .I(N__28291));
    LocalMux I__4841 (
            .O(N__28297),
            .I(N__28291));
    CascadeMux I__4840 (
            .O(N__28296),
            .I(N__28288));
    Span4Mux_v I__4839 (
            .O(N__28291),
            .I(N__28285));
    InMux I__4838 (
            .O(N__28288),
            .I(N__28282));
    Odrv4 I__4837 (
            .O(N__28285),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__4836 (
            .O(N__28282),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__4835 (
            .O(N__28277),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__4834 (
            .O(N__28274),
            .I(N__28270));
    CascadeMux I__4833 (
            .O(N__28273),
            .I(N__28267));
    InMux I__4832 (
            .O(N__28270),
            .I(N__28261));
    InMux I__4831 (
            .O(N__28267),
            .I(N__28261));
    InMux I__4830 (
            .O(N__28266),
            .I(N__28258));
    LocalMux I__4829 (
            .O(N__28261),
            .I(N__28255));
    LocalMux I__4828 (
            .O(N__28258),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv4 I__4827 (
            .O(N__28255),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__4826 (
            .O(N__28250),
            .I(N__28245));
    InMux I__4825 (
            .O(N__28249),
            .I(N__28240));
    InMux I__4824 (
            .O(N__28248),
            .I(N__28240));
    LocalMux I__4823 (
            .O(N__28245),
            .I(N__28237));
    LocalMux I__4822 (
            .O(N__28240),
            .I(N__28234));
    Span4Mux_v I__4821 (
            .O(N__28237),
            .I(N__28230));
    Sp12to4 I__4820 (
            .O(N__28234),
            .I(N__28227));
    InMux I__4819 (
            .O(N__28233),
            .I(N__28224));
    Odrv4 I__4818 (
            .O(N__28230),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv12 I__4817 (
            .O(N__28227),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__4816 (
            .O(N__28224),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__4815 (
            .O(N__28217),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__4814 (
            .O(N__28214),
            .I(N__28210));
    CascadeMux I__4813 (
            .O(N__28213),
            .I(N__28207));
    InMux I__4812 (
            .O(N__28210),
            .I(N__28201));
    InMux I__4811 (
            .O(N__28207),
            .I(N__28201));
    InMux I__4810 (
            .O(N__28206),
            .I(N__28198));
    LocalMux I__4809 (
            .O(N__28201),
            .I(N__28195));
    LocalMux I__4808 (
            .O(N__28198),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__4807 (
            .O(N__28195),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__4806 (
            .O(N__28190),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__4805 (
            .O(N__28187),
            .I(N__28184));
    InMux I__4804 (
            .O(N__28184),
            .I(N__28180));
    InMux I__4803 (
            .O(N__28183),
            .I(N__28177));
    LocalMux I__4802 (
            .O(N__28180),
            .I(N__28171));
    LocalMux I__4801 (
            .O(N__28177),
            .I(N__28171));
    InMux I__4800 (
            .O(N__28176),
            .I(N__28168));
    Span4Mux_h I__4799 (
            .O(N__28171),
            .I(N__28165));
    LocalMux I__4798 (
            .O(N__28168),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__4797 (
            .O(N__28165),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__4796 (
            .O(N__28160),
            .I(N__28157));
    LocalMux I__4795 (
            .O(N__28157),
            .I(N__28151));
    InMux I__4794 (
            .O(N__28156),
            .I(N__28144));
    InMux I__4793 (
            .O(N__28155),
            .I(N__28144));
    InMux I__4792 (
            .O(N__28154),
            .I(N__28144));
    Span4Mux_v I__4791 (
            .O(N__28151),
            .I(N__28139));
    LocalMux I__4790 (
            .O(N__28144),
            .I(N__28139));
    Odrv4 I__4789 (
            .O(N__28139),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__4788 (
            .O(N__28136),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__4787 (
            .O(N__28133),
            .I(N__28127));
    InMux I__4786 (
            .O(N__28132),
            .I(N__28127));
    LocalMux I__4785 (
            .O(N__28127),
            .I(N__28123));
    InMux I__4784 (
            .O(N__28126),
            .I(N__28120));
    Span4Mux_h I__4783 (
            .O(N__28123),
            .I(N__28117));
    LocalMux I__4782 (
            .O(N__28120),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__4781 (
            .O(N__28117),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__4780 (
            .O(N__28112),
            .I(N__28108));
    CascadeMux I__4779 (
            .O(N__28111),
            .I(N__28103));
    LocalMux I__4778 (
            .O(N__28108),
            .I(N__28100));
    InMux I__4777 (
            .O(N__28107),
            .I(N__28093));
    InMux I__4776 (
            .O(N__28106),
            .I(N__28093));
    InMux I__4775 (
            .O(N__28103),
            .I(N__28093));
    Span4Mux_h I__4774 (
            .O(N__28100),
            .I(N__28088));
    LocalMux I__4773 (
            .O(N__28093),
            .I(N__28088));
    Odrv4 I__4772 (
            .O(N__28088),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__4771 (
            .O(N__28085),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__4770 (
            .O(N__28082),
            .I(N__28079));
    InMux I__4769 (
            .O(N__28079),
            .I(N__28075));
    InMux I__4768 (
            .O(N__28078),
            .I(N__28072));
    LocalMux I__4767 (
            .O(N__28075),
            .I(N__28068));
    LocalMux I__4766 (
            .O(N__28072),
            .I(N__28065));
    InMux I__4765 (
            .O(N__28071),
            .I(N__28062));
    Span4Mux_h I__4764 (
            .O(N__28068),
            .I(N__28059));
    Span4Mux_h I__4763 (
            .O(N__28065),
            .I(N__28056));
    LocalMux I__4762 (
            .O(N__28062),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__4761 (
            .O(N__28059),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__4760 (
            .O(N__28056),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__4759 (
            .O(N__28049),
            .I(N__28046));
    LocalMux I__4758 (
            .O(N__28046),
            .I(N__28040));
    InMux I__4757 (
            .O(N__28045),
            .I(N__28035));
    InMux I__4756 (
            .O(N__28044),
            .I(N__28035));
    InMux I__4755 (
            .O(N__28043),
            .I(N__28032));
    Span4Mux_h I__4754 (
            .O(N__28040),
            .I(N__28027));
    LocalMux I__4753 (
            .O(N__28035),
            .I(N__28027));
    LocalMux I__4752 (
            .O(N__28032),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    Odrv4 I__4751 (
            .O(N__28027),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__4750 (
            .O(N__28022),
            .I(bfn_10_13_0_));
    CascadeMux I__4749 (
            .O(N__28019),
            .I(N__28015));
    CascadeMux I__4748 (
            .O(N__28018),
            .I(N__28012));
    InMux I__4747 (
            .O(N__28015),
            .I(N__28009));
    InMux I__4746 (
            .O(N__28012),
            .I(N__28006));
    LocalMux I__4745 (
            .O(N__28009),
            .I(N__28002));
    LocalMux I__4744 (
            .O(N__28006),
            .I(N__27999));
    InMux I__4743 (
            .O(N__28005),
            .I(N__27996));
    Span4Mux_h I__4742 (
            .O(N__28002),
            .I(N__27993));
    Span4Mux_h I__4741 (
            .O(N__27999),
            .I(N__27990));
    LocalMux I__4740 (
            .O(N__27996),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__4739 (
            .O(N__27993),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__4738 (
            .O(N__27990),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__4737 (
            .O(N__27983),
            .I(N__27977));
    InMux I__4736 (
            .O(N__27982),
            .I(N__27974));
    InMux I__4735 (
            .O(N__27981),
            .I(N__27971));
    InMux I__4734 (
            .O(N__27980),
            .I(N__27968));
    LocalMux I__4733 (
            .O(N__27977),
            .I(N__27961));
    LocalMux I__4732 (
            .O(N__27974),
            .I(N__27961));
    LocalMux I__4731 (
            .O(N__27971),
            .I(N__27961));
    LocalMux I__4730 (
            .O(N__27968),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__4729 (
            .O(N__27961),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__4728 (
            .O(N__27956),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__4727 (
            .O(N__27953),
            .I(N__27946));
    InMux I__4726 (
            .O(N__27952),
            .I(N__27946));
    InMux I__4725 (
            .O(N__27951),
            .I(N__27943));
    LocalMux I__4724 (
            .O(N__27946),
            .I(N__27940));
    LocalMux I__4723 (
            .O(N__27943),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__4722 (
            .O(N__27940),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__4721 (
            .O(N__27935),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__4720 (
            .O(N__27932),
            .I(N__27926));
    InMux I__4719 (
            .O(N__27931),
            .I(N__27926));
    LocalMux I__4718 (
            .O(N__27926),
            .I(N__27922));
    InMux I__4717 (
            .O(N__27925),
            .I(N__27919));
    Span4Mux_h I__4716 (
            .O(N__27922),
            .I(N__27916));
    LocalMux I__4715 (
            .O(N__27919),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__4714 (
            .O(N__27916),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__4713 (
            .O(N__27911),
            .I(N__27906));
    InMux I__4712 (
            .O(N__27910),
            .I(N__27903));
    InMux I__4711 (
            .O(N__27909),
            .I(N__27900));
    LocalMux I__4710 (
            .O(N__27906),
            .I(N__27895));
    LocalMux I__4709 (
            .O(N__27903),
            .I(N__27895));
    LocalMux I__4708 (
            .O(N__27900),
            .I(N__27889));
    Sp12to4 I__4707 (
            .O(N__27895),
            .I(N__27889));
    InMux I__4706 (
            .O(N__27894),
            .I(N__27886));
    Odrv12 I__4705 (
            .O(N__27889),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    LocalMux I__4704 (
            .O(N__27886),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__4703 (
            .O(N__27881),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__4702 (
            .O(N__27878),
            .I(N__27874));
    CascadeMux I__4701 (
            .O(N__27877),
            .I(N__27871));
    InMux I__4700 (
            .O(N__27874),
            .I(N__27865));
    InMux I__4699 (
            .O(N__27871),
            .I(N__27865));
    InMux I__4698 (
            .O(N__27870),
            .I(N__27862));
    LocalMux I__4697 (
            .O(N__27865),
            .I(N__27859));
    LocalMux I__4696 (
            .O(N__27862),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__4695 (
            .O(N__27859),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__4694 (
            .O(N__27854),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__4693 (
            .O(N__27851),
            .I(N__27845));
    InMux I__4692 (
            .O(N__27850),
            .I(N__27845));
    LocalMux I__4691 (
            .O(N__27845),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ));
    CascadeMux I__4690 (
            .O(N__27842),
            .I(N__27839));
    InMux I__4689 (
            .O(N__27839),
            .I(N__27836));
    LocalMux I__4688 (
            .O(N__27836),
            .I(N__27833));
    Odrv4 I__4687 (
            .O(N__27833),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt28 ));
    CascadeMux I__4686 (
            .O(N__27830),
            .I(N__27827));
    InMux I__4685 (
            .O(N__27827),
            .I(N__27821));
    InMux I__4684 (
            .O(N__27826),
            .I(N__27821));
    LocalMux I__4683 (
            .O(N__27821),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ));
    InMux I__4682 (
            .O(N__27818),
            .I(N__27814));
    InMux I__4681 (
            .O(N__27817),
            .I(N__27811));
    LocalMux I__4680 (
            .O(N__27814),
            .I(N__27807));
    LocalMux I__4679 (
            .O(N__27811),
            .I(N__27804));
    InMux I__4678 (
            .O(N__27810),
            .I(N__27801));
    Span4Mux_v I__4677 (
            .O(N__27807),
            .I(N__27796));
    Span4Mux_v I__4676 (
            .O(N__27804),
            .I(N__27796));
    LocalMux I__4675 (
            .O(N__27801),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__4674 (
            .O(N__27796),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__4673 (
            .O(N__27791),
            .I(N__27786));
    InMux I__4672 (
            .O(N__27790),
            .I(N__27783));
    InMux I__4671 (
            .O(N__27789),
            .I(N__27780));
    LocalMux I__4670 (
            .O(N__27786),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    LocalMux I__4669 (
            .O(N__27783),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    LocalMux I__4668 (
            .O(N__27780),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    InMux I__4667 (
            .O(N__27773),
            .I(N__27769));
    InMux I__4666 (
            .O(N__27772),
            .I(N__27765));
    LocalMux I__4665 (
            .O(N__27769),
            .I(N__27762));
    InMux I__4664 (
            .O(N__27768),
            .I(N__27759));
    LocalMux I__4663 (
            .O(N__27765),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    Odrv4 I__4662 (
            .O(N__27762),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__4661 (
            .O(N__27759),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__4660 (
            .O(N__27752),
            .I(N__27747));
    InMux I__4659 (
            .O(N__27751),
            .I(N__27744));
    InMux I__4658 (
            .O(N__27750),
            .I(N__27741));
    LocalMux I__4657 (
            .O(N__27747),
            .I(N__27736));
    LocalMux I__4656 (
            .O(N__27744),
            .I(N__27736));
    LocalMux I__4655 (
            .O(N__27741),
            .I(N__27732));
    Span4Mux_v I__4654 (
            .O(N__27736),
            .I(N__27729));
    InMux I__4653 (
            .O(N__27735),
            .I(N__27726));
    Span4Mux_v I__4652 (
            .O(N__27732),
            .I(N__27723));
    Span4Mux_h I__4651 (
            .O(N__27729),
            .I(N__27720));
    LocalMux I__4650 (
            .O(N__27726),
            .I(N__27717));
    Odrv4 I__4649 (
            .O(N__27723),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    Odrv4 I__4648 (
            .O(N__27720),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    Odrv12 I__4647 (
            .O(N__27717),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    CascadeMux I__4646 (
            .O(N__27710),
            .I(N__27707));
    InMux I__4645 (
            .O(N__27707),
            .I(N__27704));
    LocalMux I__4644 (
            .O(N__27704),
            .I(N__27699));
    InMux I__4643 (
            .O(N__27703),
            .I(N__27696));
    InMux I__4642 (
            .O(N__27702),
            .I(N__27693));
    Span4Mux_h I__4641 (
            .O(N__27699),
            .I(N__27690));
    LocalMux I__4640 (
            .O(N__27696),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__4639 (
            .O(N__27693),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    Odrv4 I__4638 (
            .O(N__27690),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__4637 (
            .O(N__27683),
            .I(N__27678));
    InMux I__4636 (
            .O(N__27682),
            .I(N__27674));
    InMux I__4635 (
            .O(N__27681),
            .I(N__27671));
    LocalMux I__4634 (
            .O(N__27678),
            .I(N__27668));
    CascadeMux I__4633 (
            .O(N__27677),
            .I(N__27665));
    LocalMux I__4632 (
            .O(N__27674),
            .I(N__27662));
    LocalMux I__4631 (
            .O(N__27671),
            .I(N__27659));
    Span4Mux_v I__4630 (
            .O(N__27668),
            .I(N__27656));
    InMux I__4629 (
            .O(N__27665),
            .I(N__27653));
    Span4Mux_h I__4628 (
            .O(N__27662),
            .I(N__27648));
    Span4Mux_v I__4627 (
            .O(N__27659),
            .I(N__27648));
    Span4Mux_h I__4626 (
            .O(N__27656),
            .I(N__27645));
    LocalMux I__4625 (
            .O(N__27653),
            .I(N__27642));
    Odrv4 I__4624 (
            .O(N__27648),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__4623 (
            .O(N__27645),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv12 I__4622 (
            .O(N__27642),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__4621 (
            .O(N__27635),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__4620 (
            .O(N__27632),
            .I(N__27628));
    InMux I__4619 (
            .O(N__27631),
            .I(N__27624));
    InMux I__4618 (
            .O(N__27628),
            .I(N__27621));
    InMux I__4617 (
            .O(N__27627),
            .I(N__27618));
    LocalMux I__4616 (
            .O(N__27624),
            .I(N__27613));
    LocalMux I__4615 (
            .O(N__27621),
            .I(N__27613));
    LocalMux I__4614 (
            .O(N__27618),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv4 I__4613 (
            .O(N__27613),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__4612 (
            .O(N__27608),
            .I(N__27601));
    InMux I__4611 (
            .O(N__27607),
            .I(N__27601));
    InMux I__4610 (
            .O(N__27606),
            .I(N__27598));
    LocalMux I__4609 (
            .O(N__27601),
            .I(N__27594));
    LocalMux I__4608 (
            .O(N__27598),
            .I(N__27591));
    InMux I__4607 (
            .O(N__27597),
            .I(N__27588));
    Span4Mux_h I__4606 (
            .O(N__27594),
            .I(N__27585));
    Span4Mux_v I__4605 (
            .O(N__27591),
            .I(N__27580));
    LocalMux I__4604 (
            .O(N__27588),
            .I(N__27580));
    Odrv4 I__4603 (
            .O(N__27585),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__4602 (
            .O(N__27580),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__4601 (
            .O(N__27575),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__4600 (
            .O(N__27572),
            .I(N__27565));
    InMux I__4599 (
            .O(N__27571),
            .I(N__27565));
    InMux I__4598 (
            .O(N__27570),
            .I(N__27562));
    LocalMux I__4597 (
            .O(N__27565),
            .I(N__27559));
    LocalMux I__4596 (
            .O(N__27562),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__4595 (
            .O(N__27559),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__4594 (
            .O(N__27554),
            .I(N__27551));
    LocalMux I__4593 (
            .O(N__27551),
            .I(N__27545));
    InMux I__4592 (
            .O(N__27550),
            .I(N__27542));
    InMux I__4591 (
            .O(N__27549),
            .I(N__27539));
    InMux I__4590 (
            .O(N__27548),
            .I(N__27536));
    Span4Mux_v I__4589 (
            .O(N__27545),
            .I(N__27531));
    LocalMux I__4588 (
            .O(N__27542),
            .I(N__27531));
    LocalMux I__4587 (
            .O(N__27539),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    LocalMux I__4586 (
            .O(N__27536),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    Odrv4 I__4585 (
            .O(N__27531),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__4584 (
            .O(N__27524),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__4583 (
            .O(N__27521),
            .I(N__27517));
    CascadeMux I__4582 (
            .O(N__27520),
            .I(N__27514));
    InMux I__4581 (
            .O(N__27517),
            .I(N__27508));
    InMux I__4580 (
            .O(N__27514),
            .I(N__27508));
    InMux I__4579 (
            .O(N__27513),
            .I(N__27505));
    LocalMux I__4578 (
            .O(N__27508),
            .I(N__27502));
    LocalMux I__4577 (
            .O(N__27505),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__4576 (
            .O(N__27502),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__4575 (
            .O(N__27497),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__4574 (
            .O(N__27494),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ));
    CascadeMux I__4573 (
            .O(N__27491),
            .I(N__27488));
    InMux I__4572 (
            .O(N__27488),
            .I(N__27485));
    LocalMux I__4571 (
            .O(N__27485),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt24 ));
    InMux I__4570 (
            .O(N__27482),
            .I(N__27476));
    InMux I__4569 (
            .O(N__27481),
            .I(N__27476));
    LocalMux I__4568 (
            .O(N__27476),
            .I(N__27473));
    Odrv12 I__4567 (
            .O(N__27473),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ));
    CascadeMux I__4566 (
            .O(N__27470),
            .I(N__27466));
    InMux I__4565 (
            .O(N__27469),
            .I(N__27461));
    InMux I__4564 (
            .O(N__27466),
            .I(N__27461));
    LocalMux I__4563 (
            .O(N__27461),
            .I(N__27458));
    Odrv12 I__4562 (
            .O(N__27458),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ));
    InMux I__4561 (
            .O(N__27455),
            .I(N__27452));
    LocalMux I__4560 (
            .O(N__27452),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ));
    InMux I__4559 (
            .O(N__27449),
            .I(N__27446));
    LocalMux I__4558 (
            .O(N__27446),
            .I(N__27442));
    InMux I__4557 (
            .O(N__27445),
            .I(N__27438));
    Span4Mux_h I__4556 (
            .O(N__27442),
            .I(N__27435));
    InMux I__4555 (
            .O(N__27441),
            .I(N__27432));
    LocalMux I__4554 (
            .O(N__27438),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    Odrv4 I__4553 (
            .O(N__27435),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    LocalMux I__4552 (
            .O(N__27432),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    InMux I__4551 (
            .O(N__27425),
            .I(N__27422));
    LocalMux I__4550 (
            .O(N__27422),
            .I(N__27419));
    Odrv4 I__4549 (
            .O(N__27419),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__4548 (
            .O(N__27416),
            .I(N__27413));
    LocalMux I__4547 (
            .O(N__27413),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ));
    CascadeMux I__4546 (
            .O(N__27410),
            .I(N__27407));
    InMux I__4545 (
            .O(N__27407),
            .I(N__27404));
    LocalMux I__4544 (
            .O(N__27404),
            .I(N__27401));
    Odrv4 I__4543 (
            .O(N__27401),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt26 ));
    InMux I__4542 (
            .O(N__27398),
            .I(N__27395));
    LocalMux I__4541 (
            .O(N__27395),
            .I(N__27392));
    Span4Mux_h I__4540 (
            .O(N__27392),
            .I(N__27388));
    InMux I__4539 (
            .O(N__27391),
            .I(N__27385));
    Odrv4 I__4538 (
            .O(N__27388),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    LocalMux I__4537 (
            .O(N__27385),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    InMux I__4536 (
            .O(N__27380),
            .I(N__27376));
    InMux I__4535 (
            .O(N__27379),
            .I(N__27373));
    LocalMux I__4534 (
            .O(N__27376),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    LocalMux I__4533 (
            .O(N__27373),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    InMux I__4532 (
            .O(N__27368),
            .I(N__27365));
    LocalMux I__4531 (
            .O(N__27365),
            .I(N__27362));
    Odrv4 I__4530 (
            .O(N__27362),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ));
    InMux I__4529 (
            .O(N__27359),
            .I(N__27356));
    LocalMux I__4528 (
            .O(N__27356),
            .I(N__27353));
    Odrv4 I__4527 (
            .O(N__27353),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    CascadeMux I__4526 (
            .O(N__27350),
            .I(N__27347));
    InMux I__4525 (
            .O(N__27347),
            .I(N__27344));
    LocalMux I__4524 (
            .O(N__27344),
            .I(N__27341));
    Span4Mux_h I__4523 (
            .O(N__27341),
            .I(N__27338));
    Odrv4 I__4522 (
            .O(N__27338),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    InMux I__4521 (
            .O(N__27335),
            .I(N__27332));
    LocalMux I__4520 (
            .O(N__27332),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ));
    CascadeMux I__4519 (
            .O(N__27329),
            .I(N__27326));
    InMux I__4518 (
            .O(N__27326),
            .I(N__27323));
    LocalMux I__4517 (
            .O(N__27323),
            .I(N__27320));
    Odrv4 I__4516 (
            .O(N__27320),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt22 ));
    InMux I__4515 (
            .O(N__27317),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ));
    InMux I__4514 (
            .O(N__27314),
            .I(N__27311));
    LocalMux I__4513 (
            .O(N__27311),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__4512 (
            .O(N__27308),
            .I(N__27305));
    LocalMux I__4511 (
            .O(N__27305),
            .I(N__27302));
    Odrv4 I__4510 (
            .O(N__27302),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    CascadeMux I__4509 (
            .O(N__27299),
            .I(N__27296));
    InMux I__4508 (
            .O(N__27296),
            .I(N__27293));
    LocalMux I__4507 (
            .O(N__27293),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__4506 (
            .O(N__27290),
            .I(N__27287));
    LocalMux I__4505 (
            .O(N__27287),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    CascadeMux I__4504 (
            .O(N__27284),
            .I(N__27281));
    InMux I__4503 (
            .O(N__27281),
            .I(N__27278));
    LocalMux I__4502 (
            .O(N__27278),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    CascadeMux I__4501 (
            .O(N__27275),
            .I(N__27272));
    InMux I__4500 (
            .O(N__27272),
            .I(N__27269));
    LocalMux I__4499 (
            .O(N__27269),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    InMux I__4498 (
            .O(N__27266),
            .I(N__27263));
    LocalMux I__4497 (
            .O(N__27263),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    CascadeMux I__4496 (
            .O(N__27260),
            .I(N__27257));
    InMux I__4495 (
            .O(N__27257),
            .I(N__27254));
    LocalMux I__4494 (
            .O(N__27254),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    CascadeMux I__4493 (
            .O(N__27251),
            .I(N__27248));
    InMux I__4492 (
            .O(N__27248),
            .I(N__27245));
    LocalMux I__4491 (
            .O(N__27245),
            .I(N__27242));
    Odrv4 I__4490 (
            .O(N__27242),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__4489 (
            .O(N__27239),
            .I(N__27236));
    LocalMux I__4488 (
            .O(N__27236),
            .I(N__27233));
    Odrv4 I__4487 (
            .O(N__27233),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__4486 (
            .O(N__27230),
            .I(N__27227));
    InMux I__4485 (
            .O(N__27227),
            .I(N__27224));
    LocalMux I__4484 (
            .O(N__27224),
            .I(N__27221));
    Odrv4 I__4483 (
            .O(N__27221),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    CascadeMux I__4482 (
            .O(N__27218),
            .I(N__27215));
    InMux I__4481 (
            .O(N__27215),
            .I(N__27212));
    LocalMux I__4480 (
            .O(N__27212),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__4479 (
            .O(N__27209),
            .I(N__27204));
    InMux I__4478 (
            .O(N__27208),
            .I(N__27201));
    InMux I__4477 (
            .O(N__27207),
            .I(N__27198));
    LocalMux I__4476 (
            .O(N__27204),
            .I(N__27195));
    LocalMux I__4475 (
            .O(N__27201),
            .I(N__27192));
    LocalMux I__4474 (
            .O(N__27198),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv12 I__4473 (
            .O(N__27195),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    Odrv4 I__4472 (
            .O(N__27192),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    CascadeMux I__4471 (
            .O(N__27185),
            .I(N__27182));
    InMux I__4470 (
            .O(N__27182),
            .I(N__27179));
    LocalMux I__4469 (
            .O(N__27179),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    InMux I__4468 (
            .O(N__27176),
            .I(N__27173));
    LocalMux I__4467 (
            .O(N__27173),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__4466 (
            .O(N__27170),
            .I(N__27167));
    LocalMux I__4465 (
            .O(N__27167),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__4464 (
            .O(N__27164),
            .I(N__27161));
    InMux I__4463 (
            .O(N__27161),
            .I(N__27158));
    LocalMux I__4462 (
            .O(N__27158),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    InMux I__4461 (
            .O(N__27155),
            .I(N__27152));
    LocalMux I__4460 (
            .O(N__27152),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__4459 (
            .O(N__27149),
            .I(N__27146));
    InMux I__4458 (
            .O(N__27146),
            .I(N__27143));
    LocalMux I__4457 (
            .O(N__27143),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__4456 (
            .O(N__27140),
            .I(N__27137));
    LocalMux I__4455 (
            .O(N__27137),
            .I(N__27134));
    Odrv4 I__4454 (
            .O(N__27134),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    CascadeMux I__4453 (
            .O(N__27131),
            .I(N__27128));
    InMux I__4452 (
            .O(N__27128),
            .I(N__27125));
    LocalMux I__4451 (
            .O(N__27125),
            .I(N__27122));
    Odrv4 I__4450 (
            .O(N__27122),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__4449 (
            .O(N__27119),
            .I(N__27116));
    LocalMux I__4448 (
            .O(N__27116),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__4447 (
            .O(N__27113),
            .I(N__27110));
    InMux I__4446 (
            .O(N__27110),
            .I(N__27107));
    LocalMux I__4445 (
            .O(N__27107),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    InMux I__4444 (
            .O(N__27104),
            .I(N__27101));
    LocalMux I__4443 (
            .O(N__27101),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    CascadeMux I__4442 (
            .O(N__27098),
            .I(N__27095));
    InMux I__4441 (
            .O(N__27095),
            .I(N__27092));
    LocalMux I__4440 (
            .O(N__27092),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__4439 (
            .O(N__27089),
            .I(N__27086));
    InMux I__4438 (
            .O(N__27086),
            .I(N__27083));
    LocalMux I__4437 (
            .O(N__27083),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__4436 (
            .O(N__27080),
            .I(N__27076));
    InMux I__4435 (
            .O(N__27079),
            .I(N__27072));
    LocalMux I__4434 (
            .O(N__27076),
            .I(N__27069));
    InMux I__4433 (
            .O(N__27075),
            .I(N__27066));
    LocalMux I__4432 (
            .O(N__27072),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    Odrv4 I__4431 (
            .O(N__27069),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    LocalMux I__4430 (
            .O(N__27066),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    CascadeMux I__4429 (
            .O(N__27059),
            .I(N__27055));
    CascadeMux I__4428 (
            .O(N__27058),
            .I(N__27052));
    InMux I__4427 (
            .O(N__27055),
            .I(N__27047));
    InMux I__4426 (
            .O(N__27052),
            .I(N__27047));
    LocalMux I__4425 (
            .O(N__27047),
            .I(N__27044));
    Odrv4 I__4424 (
            .O(N__27044),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__4423 (
            .O(N__27041),
            .I(N__27038));
    InMux I__4422 (
            .O(N__27038),
            .I(N__27035));
    LocalMux I__4421 (
            .O(N__27035),
            .I(N__27032));
    Span4Mux_v I__4420 (
            .O(N__27032),
            .I(N__27029));
    Span4Mux_v I__4419 (
            .O(N__27029),
            .I(N__27026));
    Odrv4 I__4418 (
            .O(N__27026),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__4417 (
            .O(N__27023),
            .I(N__27020));
    LocalMux I__4416 (
            .O(N__27020),
            .I(N__27016));
    InMux I__4415 (
            .O(N__27019),
            .I(N__27013));
    Span4Mux_h I__4414 (
            .O(N__27016),
            .I(N__27010));
    LocalMux I__4413 (
            .O(N__27013),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    Odrv4 I__4412 (
            .O(N__27010),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    InMux I__4411 (
            .O(N__27005),
            .I(N__27001));
    InMux I__4410 (
            .O(N__27004),
            .I(N__26998));
    LocalMux I__4409 (
            .O(N__27001),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    LocalMux I__4408 (
            .O(N__26998),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    InMux I__4407 (
            .O(N__26993),
            .I(N__26987));
    InMux I__4406 (
            .O(N__26992),
            .I(N__26987));
    LocalMux I__4405 (
            .O(N__26987),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    InMux I__4404 (
            .O(N__26984),
            .I(N__26981));
    LocalMux I__4403 (
            .O(N__26981),
            .I(N__26977));
    InMux I__4402 (
            .O(N__26980),
            .I(N__26973));
    Span4Mux_h I__4401 (
            .O(N__26977),
            .I(N__26970));
    InMux I__4400 (
            .O(N__26976),
            .I(N__26967));
    LocalMux I__4399 (
            .O(N__26973),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__4398 (
            .O(N__26970),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    LocalMux I__4397 (
            .O(N__26967),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__4396 (
            .O(N__26960),
            .I(N__26955));
    InMux I__4395 (
            .O(N__26959),
            .I(N__26952));
    InMux I__4394 (
            .O(N__26958),
            .I(N__26949));
    LocalMux I__4393 (
            .O(N__26955),
            .I(N__26946));
    LocalMux I__4392 (
            .O(N__26952),
            .I(N__26942));
    LocalMux I__4391 (
            .O(N__26949),
            .I(N__26937));
    Span4Mux_h I__4390 (
            .O(N__26946),
            .I(N__26937));
    InMux I__4389 (
            .O(N__26945),
            .I(N__26934));
    Span12Mux_v I__4388 (
            .O(N__26942),
            .I(N__26931));
    Span4Mux_v I__4387 (
            .O(N__26937),
            .I(N__26926));
    LocalMux I__4386 (
            .O(N__26934),
            .I(N__26926));
    Odrv12 I__4385 (
            .O(N__26931),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    Odrv4 I__4384 (
            .O(N__26926),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    InMux I__4383 (
            .O(N__26921),
            .I(N__26918));
    LocalMux I__4382 (
            .O(N__26918),
            .I(N__26914));
    InMux I__4381 (
            .O(N__26917),
            .I(N__26910));
    Span4Mux_v I__4380 (
            .O(N__26914),
            .I(N__26907));
    InMux I__4379 (
            .O(N__26913),
            .I(N__26904));
    LocalMux I__4378 (
            .O(N__26910),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    Odrv4 I__4377 (
            .O(N__26907),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    LocalMux I__4376 (
            .O(N__26904),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    InMux I__4375 (
            .O(N__26897),
            .I(N__26892));
    InMux I__4374 (
            .O(N__26896),
            .I(N__26889));
    InMux I__4373 (
            .O(N__26895),
            .I(N__26886));
    LocalMux I__4372 (
            .O(N__26892),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    LocalMux I__4371 (
            .O(N__26889),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    LocalMux I__4370 (
            .O(N__26886),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    InMux I__4369 (
            .O(N__26879),
            .I(N__26876));
    LocalMux I__4368 (
            .O(N__26876),
            .I(N__26873));
    Span4Mux_h I__4367 (
            .O(N__26873),
            .I(N__26868));
    InMux I__4366 (
            .O(N__26872),
            .I(N__26865));
    InMux I__4365 (
            .O(N__26871),
            .I(N__26862));
    Span4Mux_v I__4364 (
            .O(N__26868),
            .I(N__26859));
    LocalMux I__4363 (
            .O(N__26865),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    LocalMux I__4362 (
            .O(N__26862),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    Odrv4 I__4361 (
            .O(N__26859),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    InMux I__4360 (
            .O(N__26852),
            .I(N__26848));
    InMux I__4359 (
            .O(N__26851),
            .I(N__26844));
    LocalMux I__4358 (
            .O(N__26848),
            .I(N__26841));
    InMux I__4357 (
            .O(N__26847),
            .I(N__26838));
    LocalMux I__4356 (
            .O(N__26844),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    Odrv4 I__4355 (
            .O(N__26841),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    LocalMux I__4354 (
            .O(N__26838),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    InMux I__4353 (
            .O(N__26831),
            .I(N__26828));
    LocalMux I__4352 (
            .O(N__26828),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__4351 (
            .O(N__26825),
            .I(N__26822));
    InMux I__4350 (
            .O(N__26822),
            .I(N__26819));
    LocalMux I__4349 (
            .O(N__26819),
            .I(N__26816));
    Odrv4 I__4348 (
            .O(N__26816),
            .I(\pwm_generator_inst.threshold_5 ));
    InMux I__4347 (
            .O(N__26813),
            .I(N__26810));
    LocalMux I__4346 (
            .O(N__26810),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__4345 (
            .O(N__26807),
            .I(N__26804));
    InMux I__4344 (
            .O(N__26804),
            .I(N__26801));
    LocalMux I__4343 (
            .O(N__26801),
            .I(N__26798));
    Span4Mux_h I__4342 (
            .O(N__26798),
            .I(N__26795));
    Odrv4 I__4341 (
            .O(N__26795),
            .I(\pwm_generator_inst.un14_counter_6 ));
    InMux I__4340 (
            .O(N__26792),
            .I(N__26789));
    LocalMux I__4339 (
            .O(N__26789),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__4338 (
            .O(N__26786),
            .I(N__26783));
    InMux I__4337 (
            .O(N__26783),
            .I(N__26780));
    LocalMux I__4336 (
            .O(N__26780),
            .I(\pwm_generator_inst.un14_counter_7 ));
    InMux I__4335 (
            .O(N__26777),
            .I(N__26774));
    LocalMux I__4334 (
            .O(N__26774),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__4333 (
            .O(N__26771),
            .I(N__26768));
    InMux I__4332 (
            .O(N__26768),
            .I(N__26765));
    LocalMux I__4331 (
            .O(N__26765),
            .I(N__26762));
    Odrv4 I__4330 (
            .O(N__26762),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__4329 (
            .O(N__26759),
            .I(N__26756));
    LocalMux I__4328 (
            .O(N__26756),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__4327 (
            .O(N__26753),
            .I(N__26750));
    InMux I__4326 (
            .O(N__26750),
            .I(N__26747));
    LocalMux I__4325 (
            .O(N__26747),
            .I(\pwm_generator_inst.threshold_9 ));
    InMux I__4324 (
            .O(N__26744),
            .I(N__26741));
    LocalMux I__4323 (
            .O(N__26741),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__4322 (
            .O(N__26738),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__4321 (
            .O(N__26735),
            .I(N__26732));
    LocalMux I__4320 (
            .O(N__26732),
            .I(N__26729));
    Span4Mux_s2_v I__4319 (
            .O(N__26729),
            .I(N__26726));
    Sp12to4 I__4318 (
            .O(N__26726),
            .I(N__26723));
    Span12Mux_h I__4317 (
            .O(N__26723),
            .I(N__26720));
    Span12Mux_v I__4316 (
            .O(N__26720),
            .I(N__26717));
    Odrv12 I__4315 (
            .O(N__26717),
            .I(pwm_output_c));
    IoInMux I__4314 (
            .O(N__26714),
            .I(N__26711));
    LocalMux I__4313 (
            .O(N__26711),
            .I(s3_phy_c));
    InMux I__4312 (
            .O(N__26708),
            .I(N__26705));
    LocalMux I__4311 (
            .O(N__26705),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__4310 (
            .O(N__26702),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__4309 (
            .O(N__26699),
            .I(N__26696));
    LocalMux I__4308 (
            .O(N__26696),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__4307 (
            .O(N__26693),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__4306 (
            .O(N__26690),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__4305 (
            .O(N__26687),
            .I(N__26683));
    InMux I__4304 (
            .O(N__26686),
            .I(N__26680));
    LocalMux I__4303 (
            .O(N__26683),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__4302 (
            .O(N__26680),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__4301 (
            .O(N__26675),
            .I(N__26672));
    LocalMux I__4300 (
            .O(N__26672),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    CascadeMux I__4299 (
            .O(N__26669),
            .I(N__26666));
    InMux I__4298 (
            .O(N__26666),
            .I(N__26663));
    LocalMux I__4297 (
            .O(N__26663),
            .I(N__26660));
    Odrv4 I__4296 (
            .O(N__26660),
            .I(\pwm_generator_inst.threshold_0 ));
    InMux I__4295 (
            .O(N__26657),
            .I(N__26654));
    LocalMux I__4294 (
            .O(N__26654),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__4293 (
            .O(N__26651),
            .I(N__26648));
    InMux I__4292 (
            .O(N__26648),
            .I(N__26645));
    LocalMux I__4291 (
            .O(N__26645),
            .I(\pwm_generator_inst.un14_counter_1 ));
    InMux I__4290 (
            .O(N__26642),
            .I(N__26639));
    LocalMux I__4289 (
            .O(N__26639),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__4288 (
            .O(N__26636),
            .I(N__26633));
    InMux I__4287 (
            .O(N__26633),
            .I(N__26630));
    LocalMux I__4286 (
            .O(N__26630),
            .I(\pwm_generator_inst.threshold_2 ));
    InMux I__4285 (
            .O(N__26627),
            .I(N__26624));
    LocalMux I__4284 (
            .O(N__26624),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__4283 (
            .O(N__26621),
            .I(N__26618));
    InMux I__4282 (
            .O(N__26618),
            .I(N__26615));
    LocalMux I__4281 (
            .O(N__26615),
            .I(\pwm_generator_inst.threshold_3 ));
    InMux I__4280 (
            .O(N__26612),
            .I(N__26609));
    LocalMux I__4279 (
            .O(N__26609),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__4278 (
            .O(N__26606),
            .I(N__26603));
    InMux I__4277 (
            .O(N__26603),
            .I(N__26600));
    LocalMux I__4276 (
            .O(N__26600),
            .I(N__26597));
    Odrv4 I__4275 (
            .O(N__26597),
            .I(\pwm_generator_inst.threshold_4 ));
    InMux I__4274 (
            .O(N__26594),
            .I(N__26591));
    LocalMux I__4273 (
            .O(N__26591),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__4272 (
            .O(N__26588),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__4271 (
            .O(N__26585),
            .I(N__26582));
    LocalMux I__4270 (
            .O(N__26582),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__4269 (
            .O(N__26579),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__4268 (
            .O(N__26576),
            .I(N__26573));
    LocalMux I__4267 (
            .O(N__26573),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__4266 (
            .O(N__26570),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__4265 (
            .O(N__26567),
            .I(N__26564));
    LocalMux I__4264 (
            .O(N__26564),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__4263 (
            .O(N__26561),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__4262 (
            .O(N__26558),
            .I(N__26555));
    LocalMux I__4261 (
            .O(N__26555),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__4260 (
            .O(N__26552),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__4259 (
            .O(N__26549),
            .I(N__26546));
    LocalMux I__4258 (
            .O(N__26546),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__4257 (
            .O(N__26543),
            .I(bfn_9_20_0_));
    InMux I__4256 (
            .O(N__26540),
            .I(N__26537));
    LocalMux I__4255 (
            .O(N__26537),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__4254 (
            .O(N__26534),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__4253 (
            .O(N__26531),
            .I(N__26528));
    LocalMux I__4252 (
            .O(N__26528),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__4251 (
            .O(N__26525),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__4250 (
            .O(N__26522),
            .I(bfn_9_18_0_));
    InMux I__4249 (
            .O(N__26519),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__4248 (
            .O(N__26516),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__4247 (
            .O(N__26513),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__4246 (
            .O(N__26510),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__4245 (
            .O(N__26507),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__4244 (
            .O(N__26504),
            .I(N__26501));
    LocalMux I__4243 (
            .O(N__26501),
            .I(\current_shift_inst.control_input_18 ));
    InMux I__4242 (
            .O(N__26498),
            .I(N__26495));
    LocalMux I__4241 (
            .O(N__26495),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__4240 (
            .O(N__26492),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__4239 (
            .O(N__26489),
            .I(N__26486));
    LocalMux I__4238 (
            .O(N__26486),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__4237 (
            .O(N__26483),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__4236 (
            .O(N__26480),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__4235 (
            .O(N__26477),
            .I(bfn_9_17_0_));
    InMux I__4234 (
            .O(N__26474),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__4233 (
            .O(N__26471),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__4232 (
            .O(N__26468),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__4231 (
            .O(N__26465),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__4230 (
            .O(N__26462),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__4229 (
            .O(N__26459),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__4228 (
            .O(N__26456),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__4227 (
            .O(N__26453),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__4226 (
            .O(N__26450),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__4225 (
            .O(N__26447),
            .I(bfn_9_16_0_));
    InMux I__4224 (
            .O(N__26444),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__4223 (
            .O(N__26441),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__4222 (
            .O(N__26438),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__4221 (
            .O(N__26435),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__4220 (
            .O(N__26432),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__4219 (
            .O(N__26429),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__4218 (
            .O(N__26426),
            .I(N__26423));
    LocalMux I__4217 (
            .O(N__26423),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ));
    InMux I__4216 (
            .O(N__26420),
            .I(N__26417));
    LocalMux I__4215 (
            .O(N__26417),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    InMux I__4214 (
            .O(N__26414),
            .I(bfn_9_15_0_));
    InMux I__4213 (
            .O(N__26411),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__4212 (
            .O(N__26408),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__4211 (
            .O(N__26405),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__4210 (
            .O(N__26402),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__4209 (
            .O(N__26399),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__4208 (
            .O(N__26396),
            .I(N__26393));
    LocalMux I__4207 (
            .O(N__26393),
            .I(N__26390));
    Odrv4 I__4206 (
            .O(N__26390),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ));
    InMux I__4205 (
            .O(N__26387),
            .I(N__26384));
    LocalMux I__4204 (
            .O(N__26384),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    CascadeMux I__4203 (
            .O(N__26381),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_ ));
    InMux I__4202 (
            .O(N__26378),
            .I(N__26375));
    LocalMux I__4201 (
            .O(N__26375),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ));
    CascadeMux I__4200 (
            .O(N__26372),
            .I(N__26369));
    InMux I__4199 (
            .O(N__26369),
            .I(N__26366));
    LocalMux I__4198 (
            .O(N__26366),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    InMux I__4197 (
            .O(N__26363),
            .I(N__26360));
    LocalMux I__4196 (
            .O(N__26360),
            .I(N__26355));
    InMux I__4195 (
            .O(N__26359),
            .I(N__26352));
    InMux I__4194 (
            .O(N__26358),
            .I(N__26349));
    Span4Mux_h I__4193 (
            .O(N__26355),
            .I(N__26344));
    LocalMux I__4192 (
            .O(N__26352),
            .I(N__26344));
    LocalMux I__4191 (
            .O(N__26349),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv4 I__4190 (
            .O(N__26344),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    InMux I__4189 (
            .O(N__26339),
            .I(N__26336));
    LocalMux I__4188 (
            .O(N__26336),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__4187 (
            .O(N__26333),
            .I(N__26324));
    InMux I__4186 (
            .O(N__26332),
            .I(N__26324));
    InMux I__4185 (
            .O(N__26331),
            .I(N__26324));
    LocalMux I__4184 (
            .O(N__26324),
            .I(N__26321));
    Span4Mux_h I__4183 (
            .O(N__26321),
            .I(N__26318));
    Odrv4 I__4182 (
            .O(N__26318),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    InMux I__4181 (
            .O(N__26315),
            .I(N__26312));
    LocalMux I__4180 (
            .O(N__26312),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__4179 (
            .O(N__26309),
            .I(N__26303));
    InMux I__4178 (
            .O(N__26308),
            .I(N__26303));
    LocalMux I__4177 (
            .O(N__26303),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ));
    CascadeMux I__4176 (
            .O(N__26300),
            .I(N__26297));
    InMux I__4175 (
            .O(N__26297),
            .I(N__26294));
    LocalMux I__4174 (
            .O(N__26294),
            .I(N__26291));
    Span4Mux_v I__4173 (
            .O(N__26291),
            .I(N__26288));
    Odrv4 I__4172 (
            .O(N__26288),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    InMux I__4171 (
            .O(N__26285),
            .I(N__26282));
    LocalMux I__4170 (
            .O(N__26282),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__4169 (
            .O(N__26279),
            .I(N__26276));
    LocalMux I__4168 (
            .O(N__26276),
            .I(N__26273));
    Odrv4 I__4167 (
            .O(N__26273),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    CascadeMux I__4166 (
            .O(N__26270),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    CascadeMux I__4165 (
            .O(N__26267),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ));
    InMux I__4164 (
            .O(N__26264),
            .I(N__26260));
    InMux I__4163 (
            .O(N__26263),
            .I(N__26257));
    LocalMux I__4162 (
            .O(N__26260),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    LocalMux I__4161 (
            .O(N__26257),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    CascadeMux I__4160 (
            .O(N__26252),
            .I(elapsed_time_ns_1_RNITUBN9_0_10_cascade_));
    InMux I__4159 (
            .O(N__26249),
            .I(N__26246));
    LocalMux I__4158 (
            .O(N__26246),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__4157 (
            .O(N__26243),
            .I(N__26240));
    LocalMux I__4156 (
            .O(N__26240),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ));
    CascadeMux I__4155 (
            .O(N__26237),
            .I(elapsed_time_ns_1_RNIL73T9_0_9_cascade_));
    InMux I__4154 (
            .O(N__26234),
            .I(N__26231));
    LocalMux I__4153 (
            .O(N__26231),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__4152 (
            .O(N__26228),
            .I(N__26225));
    LocalMux I__4151 (
            .O(N__26225),
            .I(N__26222));
    Span4Mux_v I__4150 (
            .O(N__26222),
            .I(N__26219));
    Odrv4 I__4149 (
            .O(N__26219),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ));
    CascadeMux I__4148 (
            .O(N__26216),
            .I(elapsed_time_ns_1_RNI14DN9_0_23_cascade_));
    CascadeMux I__4147 (
            .O(N__26213),
            .I(N__26210));
    InMux I__4146 (
            .O(N__26210),
            .I(N__26204));
    InMux I__4145 (
            .O(N__26209),
            .I(N__26204));
    LocalMux I__4144 (
            .O(N__26204),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    CascadeMux I__4143 (
            .O(N__26201),
            .I(elapsed_time_ns_1_RNI03DN9_0_22_cascade_));
    InMux I__4142 (
            .O(N__26198),
            .I(N__26192));
    InMux I__4141 (
            .O(N__26197),
            .I(N__26192));
    LocalMux I__4140 (
            .O(N__26192),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ));
    InMux I__4139 (
            .O(N__26189),
            .I(N__26186));
    LocalMux I__4138 (
            .O(N__26186),
            .I(N__26181));
    InMux I__4137 (
            .O(N__26185),
            .I(N__26178));
    InMux I__4136 (
            .O(N__26184),
            .I(N__26175));
    Span4Mux_v I__4135 (
            .O(N__26181),
            .I(N__26170));
    LocalMux I__4134 (
            .O(N__26178),
            .I(N__26170));
    LocalMux I__4133 (
            .O(N__26175),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    Odrv4 I__4132 (
            .O(N__26170),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    InMux I__4131 (
            .O(N__26165),
            .I(N__26162));
    LocalMux I__4130 (
            .O(N__26162),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__4129 (
            .O(N__26159),
            .I(N__26155));
    InMux I__4128 (
            .O(N__26158),
            .I(N__26152));
    LocalMux I__4127 (
            .O(N__26155),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    LocalMux I__4126 (
            .O(N__26152),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    InMux I__4125 (
            .O(N__26147),
            .I(N__26141));
    InMux I__4124 (
            .O(N__26146),
            .I(N__26141));
    LocalMux I__4123 (
            .O(N__26141),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    InMux I__4122 (
            .O(N__26138),
            .I(N__26134));
    InMux I__4121 (
            .O(N__26137),
            .I(N__26131));
    LocalMux I__4120 (
            .O(N__26134),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    LocalMux I__4119 (
            .O(N__26131),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    CascadeMux I__4118 (
            .O(N__26126),
            .I(N__26123));
    InMux I__4117 (
            .O(N__26123),
            .I(N__26117));
    InMux I__4116 (
            .O(N__26122),
            .I(N__26117));
    LocalMux I__4115 (
            .O(N__26117),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    CascadeMux I__4114 (
            .O(N__26114),
            .I(N__26111));
    InMux I__4113 (
            .O(N__26111),
            .I(N__26105));
    InMux I__4112 (
            .O(N__26110),
            .I(N__26105));
    LocalMux I__4111 (
            .O(N__26105),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    InMux I__4110 (
            .O(N__26102),
            .I(N__26097));
    InMux I__4109 (
            .O(N__26101),
            .I(N__26094));
    InMux I__4108 (
            .O(N__26100),
            .I(N__26091));
    LocalMux I__4107 (
            .O(N__26097),
            .I(N__26088));
    LocalMux I__4106 (
            .O(N__26094),
            .I(N__26085));
    LocalMux I__4105 (
            .O(N__26091),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__4104 (
            .O(N__26088),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__4103 (
            .O(N__26085),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__4102 (
            .O(N__26078),
            .I(N__26074));
    InMux I__4101 (
            .O(N__26077),
            .I(N__26070));
    LocalMux I__4100 (
            .O(N__26074),
            .I(N__26067));
    InMux I__4099 (
            .O(N__26073),
            .I(N__26064));
    LocalMux I__4098 (
            .O(N__26070),
            .I(N__26061));
    Span4Mux_h I__4097 (
            .O(N__26067),
            .I(N__26053));
    LocalMux I__4096 (
            .O(N__26064),
            .I(N__26053));
    Span4Mux_h I__4095 (
            .O(N__26061),
            .I(N__26053));
    InMux I__4094 (
            .O(N__26060),
            .I(N__26050));
    Span4Mux_v I__4093 (
            .O(N__26053),
            .I(N__26045));
    LocalMux I__4092 (
            .O(N__26050),
            .I(N__26045));
    Odrv4 I__4091 (
            .O(N__26045),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__4090 (
            .O(N__26042),
            .I(N__26038));
    InMux I__4089 (
            .O(N__26041),
            .I(N__26034));
    LocalMux I__4088 (
            .O(N__26038),
            .I(N__26031));
    InMux I__4087 (
            .O(N__26037),
            .I(N__26028));
    LocalMux I__4086 (
            .O(N__26034),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv4 I__4085 (
            .O(N__26031),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    LocalMux I__4084 (
            .O(N__26028),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    InMux I__4083 (
            .O(N__26021),
            .I(N__26018));
    LocalMux I__4082 (
            .O(N__26018),
            .I(N__26015));
    Span4Mux_v I__4081 (
            .O(N__26015),
            .I(N__26011));
    InMux I__4080 (
            .O(N__26014),
            .I(N__26008));
    Odrv4 I__4079 (
            .O(N__26011),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__4078 (
            .O(N__26008),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    CascadeMux I__4077 (
            .O(N__26003),
            .I(N__26000));
    InMux I__4076 (
            .O(N__26000),
            .I(N__25997));
    LocalMux I__4075 (
            .O(N__25997),
            .I(N__25994));
    Span4Mux_v I__4074 (
            .O(N__25994),
            .I(N__25991));
    Odrv4 I__4073 (
            .O(N__25991),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt22 ));
    CascadeMux I__4072 (
            .O(N__25988),
            .I(N__25983));
    InMux I__4071 (
            .O(N__25987),
            .I(N__25980));
    InMux I__4070 (
            .O(N__25986),
            .I(N__25975));
    InMux I__4069 (
            .O(N__25983),
            .I(N__25975));
    LocalMux I__4068 (
            .O(N__25980),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    LocalMux I__4067 (
            .O(N__25975),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__4066 (
            .O(N__25970),
            .I(N__25965));
    InMux I__4065 (
            .O(N__25969),
            .I(N__25960));
    InMux I__4064 (
            .O(N__25968),
            .I(N__25960));
    LocalMux I__4063 (
            .O(N__25965),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    LocalMux I__4062 (
            .O(N__25960),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__4061 (
            .O(N__25955),
            .I(N__25950));
    InMux I__4060 (
            .O(N__25954),
            .I(N__25947));
    InMux I__4059 (
            .O(N__25953),
            .I(N__25944));
    LocalMux I__4058 (
            .O(N__25950),
            .I(N__25941));
    LocalMux I__4057 (
            .O(N__25947),
            .I(N__25938));
    LocalMux I__4056 (
            .O(N__25944),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__4055 (
            .O(N__25941),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__4054 (
            .O(N__25938),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__4053 (
            .O(N__25931),
            .I(N__25928));
    InMux I__4052 (
            .O(N__25928),
            .I(N__25923));
    InMux I__4051 (
            .O(N__25927),
            .I(N__25920));
    InMux I__4050 (
            .O(N__25926),
            .I(N__25917));
    LocalMux I__4049 (
            .O(N__25923),
            .I(N__25914));
    LocalMux I__4048 (
            .O(N__25920),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__4047 (
            .O(N__25917),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    Odrv4 I__4046 (
            .O(N__25914),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__4045 (
            .O(N__25907),
            .I(N__25904));
    InMux I__4044 (
            .O(N__25904),
            .I(N__25900));
    InMux I__4043 (
            .O(N__25903),
            .I(N__25897));
    LocalMux I__4042 (
            .O(N__25900),
            .I(N__25894));
    LocalMux I__4041 (
            .O(N__25897),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    Odrv4 I__4040 (
            .O(N__25894),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__4039 (
            .O(N__25889),
            .I(N__25885));
    InMux I__4038 (
            .O(N__25888),
            .I(N__25882));
    LocalMux I__4037 (
            .O(N__25885),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    LocalMux I__4036 (
            .O(N__25882),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__4035 (
            .O(N__25877),
            .I(N__25874));
    InMux I__4034 (
            .O(N__25874),
            .I(N__25871));
    LocalMux I__4033 (
            .O(N__25871),
            .I(N__25868));
    Sp12to4 I__4032 (
            .O(N__25868),
            .I(N__25865));
    Odrv12 I__4031 (
            .O(N__25865),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    InMux I__4030 (
            .O(N__25862),
            .I(N__25859));
    LocalMux I__4029 (
            .O(N__25859),
            .I(N__25856));
    Span4Mux_v I__4028 (
            .O(N__25856),
            .I(N__25853));
    Odrv4 I__4027 (
            .O(N__25853),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    CascadeMux I__4026 (
            .O(N__25850),
            .I(elapsed_time_ns_1_RNI57CN9_0_18_cascade_));
    InMux I__4025 (
            .O(N__25847),
            .I(N__25841));
    InMux I__4024 (
            .O(N__25846),
            .I(N__25841));
    LocalMux I__4023 (
            .O(N__25841),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    InMux I__4022 (
            .O(N__25838),
            .I(N__25833));
    InMux I__4021 (
            .O(N__25837),
            .I(N__25828));
    InMux I__4020 (
            .O(N__25836),
            .I(N__25828));
    LocalMux I__4019 (
            .O(N__25833),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__4018 (
            .O(N__25828),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__4017 (
            .O(N__25823),
            .I(N__25818));
    InMux I__4016 (
            .O(N__25822),
            .I(N__25813));
    InMux I__4015 (
            .O(N__25821),
            .I(N__25813));
    LocalMux I__4014 (
            .O(N__25818),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__4013 (
            .O(N__25813),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    CascadeMux I__4012 (
            .O(N__25808),
            .I(N__25805));
    InMux I__4011 (
            .O(N__25805),
            .I(N__25802));
    LocalMux I__4010 (
            .O(N__25802),
            .I(N__25799));
    Span4Mux_v I__4009 (
            .O(N__25799),
            .I(N__25796));
    Odrv4 I__4008 (
            .O(N__25796),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    CascadeMux I__4007 (
            .O(N__25793),
            .I(elapsed_time_ns_1_RNI24CN9_0_15_cascade_));
    InMux I__4006 (
            .O(N__25790),
            .I(N__25787));
    LocalMux I__4005 (
            .O(N__25787),
            .I(N__25784));
    Span4Mux_v I__4004 (
            .O(N__25784),
            .I(N__25781));
    Odrv4 I__4003 (
            .O(N__25781),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    CascadeMux I__4002 (
            .O(N__25778),
            .I(N__25775));
    InMux I__4001 (
            .O(N__25775),
            .I(N__25772));
    LocalMux I__4000 (
            .O(N__25772),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ));
    InMux I__3999 (
            .O(N__25769),
            .I(N__25766));
    LocalMux I__3998 (
            .O(N__25766),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ));
    InMux I__3997 (
            .O(N__25763),
            .I(N__25760));
    LocalMux I__3996 (
            .O(N__25760),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ));
    CascadeMux I__3995 (
            .O(N__25757),
            .I(N__25754));
    InMux I__3994 (
            .O(N__25754),
            .I(N__25751));
    LocalMux I__3993 (
            .O(N__25751),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ));
    InMux I__3992 (
            .O(N__25748),
            .I(N__25745));
    LocalMux I__3991 (
            .O(N__25745),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ));
    InMux I__3990 (
            .O(N__25742),
            .I(N__25739));
    LocalMux I__3989 (
            .O(N__25739),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ));
    InMux I__3988 (
            .O(N__25736),
            .I(N__25721));
    InMux I__3987 (
            .O(N__25735),
            .I(N__25721));
    InMux I__3986 (
            .O(N__25734),
            .I(N__25721));
    InMux I__3985 (
            .O(N__25733),
            .I(N__25721));
    InMux I__3984 (
            .O(N__25732),
            .I(N__25721));
    LocalMux I__3983 (
            .O(N__25721),
            .I(N__25713));
    InMux I__3982 (
            .O(N__25720),
            .I(N__25702));
    InMux I__3981 (
            .O(N__25719),
            .I(N__25702));
    InMux I__3980 (
            .O(N__25718),
            .I(N__25702));
    InMux I__3979 (
            .O(N__25717),
            .I(N__25702));
    InMux I__3978 (
            .O(N__25716),
            .I(N__25702));
    Sp12to4 I__3977 (
            .O(N__25713),
            .I(N__25697));
    LocalMux I__3976 (
            .O(N__25702),
            .I(N__25697));
    Span12Mux_s7_v I__3975 (
            .O(N__25697),
            .I(N__25694));
    Odrv12 I__3974 (
            .O(N__25694),
            .I(\pwm_generator_inst.N_17 ));
    InMux I__3973 (
            .O(N__25691),
            .I(N__25671));
    InMux I__3972 (
            .O(N__25690),
            .I(N__25671));
    InMux I__3971 (
            .O(N__25689),
            .I(N__25671));
    InMux I__3970 (
            .O(N__25688),
            .I(N__25671));
    InMux I__3969 (
            .O(N__25687),
            .I(N__25671));
    InMux I__3968 (
            .O(N__25686),
            .I(N__25660));
    InMux I__3967 (
            .O(N__25685),
            .I(N__25660));
    InMux I__3966 (
            .O(N__25684),
            .I(N__25660));
    InMux I__3965 (
            .O(N__25683),
            .I(N__25660));
    InMux I__3964 (
            .O(N__25682),
            .I(N__25660));
    LocalMux I__3963 (
            .O(N__25671),
            .I(N__25657));
    LocalMux I__3962 (
            .O(N__25660),
            .I(N__25654));
    Span4Mux_h I__3961 (
            .O(N__25657),
            .I(N__25649));
    Span4Mux_v I__3960 (
            .O(N__25654),
            .I(N__25649));
    Span4Mux_h I__3959 (
            .O(N__25649),
            .I(N__25646));
    Odrv4 I__3958 (
            .O(N__25646),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__3957 (
            .O(N__25643),
            .I(N__25640));
    InMux I__3956 (
            .O(N__25640),
            .I(N__25637));
    LocalMux I__3955 (
            .O(N__25637),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ));
    InMux I__3954 (
            .O(N__25634),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__3953 (
            .O(N__25631),
            .I(N__25628));
    LocalMux I__3952 (
            .O(N__25628),
            .I(N__25624));
    InMux I__3951 (
            .O(N__25627),
            .I(N__25621));
    Span4Mux_v I__3950 (
            .O(N__25624),
            .I(N__25618));
    LocalMux I__3949 (
            .O(N__25621),
            .I(N__25615));
    Sp12to4 I__3948 (
            .O(N__25618),
            .I(N__25612));
    Span4Mux_h I__3947 (
            .O(N__25615),
            .I(N__25609));
    Span12Mux_s8_h I__3946 (
            .O(N__25612),
            .I(N__25606));
    Odrv4 I__3945 (
            .O(N__25609),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv12 I__3944 (
            .O(N__25606),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__3943 (
            .O(N__25601),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__3942 (
            .O(N__25598),
            .I(N__25594));
    InMux I__3941 (
            .O(N__25597),
            .I(N__25591));
    LocalMux I__3940 (
            .O(N__25594),
            .I(N__25588));
    LocalMux I__3939 (
            .O(N__25591),
            .I(N__25585));
    Span12Mux_s8_h I__3938 (
            .O(N__25588),
            .I(N__25582));
    Span4Mux_v I__3937 (
            .O(N__25585),
            .I(N__25579));
    Span12Mux_v I__3936 (
            .O(N__25582),
            .I(N__25576));
    Odrv4 I__3935 (
            .O(N__25579),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv12 I__3934 (
            .O(N__25576),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__3933 (
            .O(N__25571),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__3932 (
            .O(N__25568),
            .I(N__25564));
    InMux I__3931 (
            .O(N__25567),
            .I(N__25561));
    LocalMux I__3930 (
            .O(N__25564),
            .I(N__25558));
    LocalMux I__3929 (
            .O(N__25561),
            .I(N__25555));
    Span12Mux_s7_v I__3928 (
            .O(N__25558),
            .I(N__25552));
    Span4Mux_h I__3927 (
            .O(N__25555),
            .I(N__25549));
    Span12Mux_v I__3926 (
            .O(N__25552),
            .I(N__25546));
    Odrv4 I__3925 (
            .O(N__25549),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv12 I__3924 (
            .O(N__25546),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__3923 (
            .O(N__25541),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__3922 (
            .O(N__25538),
            .I(N__25535));
    LocalMux I__3921 (
            .O(N__25535),
            .I(N__25532));
    Span4Mux_v I__3920 (
            .O(N__25532),
            .I(N__25528));
    InMux I__3919 (
            .O(N__25531),
            .I(N__25525));
    Span4Mux_v I__3918 (
            .O(N__25528),
            .I(N__25522));
    LocalMux I__3917 (
            .O(N__25525),
            .I(N__25519));
    Sp12to4 I__3916 (
            .O(N__25522),
            .I(N__25516));
    Span4Mux_h I__3915 (
            .O(N__25519),
            .I(N__25513));
    Span12Mux_s8_h I__3914 (
            .O(N__25516),
            .I(N__25510));
    Odrv4 I__3913 (
            .O(N__25513),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv12 I__3912 (
            .O(N__25510),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__3911 (
            .O(N__25505),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__3910 (
            .O(N__25502),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__3909 (
            .O(N__25499),
            .I(N__25480));
    InMux I__3908 (
            .O(N__25498),
            .I(N__25463));
    InMux I__3907 (
            .O(N__25497),
            .I(N__25463));
    InMux I__3906 (
            .O(N__25496),
            .I(N__25463));
    InMux I__3905 (
            .O(N__25495),
            .I(N__25463));
    InMux I__3904 (
            .O(N__25494),
            .I(N__25463));
    InMux I__3903 (
            .O(N__25493),
            .I(N__25463));
    InMux I__3902 (
            .O(N__25492),
            .I(N__25463));
    InMux I__3901 (
            .O(N__25491),
            .I(N__25463));
    InMux I__3900 (
            .O(N__25490),
            .I(N__25446));
    InMux I__3899 (
            .O(N__25489),
            .I(N__25446));
    InMux I__3898 (
            .O(N__25488),
            .I(N__25446));
    InMux I__3897 (
            .O(N__25487),
            .I(N__25446));
    InMux I__3896 (
            .O(N__25486),
            .I(N__25446));
    InMux I__3895 (
            .O(N__25485),
            .I(N__25446));
    InMux I__3894 (
            .O(N__25484),
            .I(N__25446));
    InMux I__3893 (
            .O(N__25483),
            .I(N__25446));
    LocalMux I__3892 (
            .O(N__25480),
            .I(N__25443));
    LocalMux I__3891 (
            .O(N__25463),
            .I(N__25435));
    LocalMux I__3890 (
            .O(N__25446),
            .I(N__25435));
    Span4Mux_v I__3889 (
            .O(N__25443),
            .I(N__25435));
    InMux I__3888 (
            .O(N__25442),
            .I(N__25432));
    Span4Mux_v I__3887 (
            .O(N__25435),
            .I(N__25429));
    LocalMux I__3886 (
            .O(N__25432),
            .I(N__25426));
    Sp12to4 I__3885 (
            .O(N__25429),
            .I(N__25423));
    Span4Mux_h I__3884 (
            .O(N__25426),
            .I(N__25420));
    Span12Mux_s8_h I__3883 (
            .O(N__25423),
            .I(N__25417));
    Odrv4 I__3882 (
            .O(N__25420),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv12 I__3881 (
            .O(N__25417),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    CascadeMux I__3880 (
            .O(N__25412),
            .I(N__25409));
    InMux I__3879 (
            .O(N__25409),
            .I(N__25406));
    LocalMux I__3878 (
            .O(N__25406),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ));
    CascadeMux I__3877 (
            .O(N__25403),
            .I(N__25400));
    InMux I__3876 (
            .O(N__25400),
            .I(N__25397));
    LocalMux I__3875 (
            .O(N__25397),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ));
    CascadeMux I__3874 (
            .O(N__25394),
            .I(N__25391));
    InMux I__3873 (
            .O(N__25391),
            .I(N__25388));
    LocalMux I__3872 (
            .O(N__25388),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ));
    InMux I__3871 (
            .O(N__25385),
            .I(N__25381));
    InMux I__3870 (
            .O(N__25384),
            .I(N__25378));
    LocalMux I__3869 (
            .O(N__25381),
            .I(N__25375));
    LocalMux I__3868 (
            .O(N__25378),
            .I(N__25372));
    Span4Mux_v I__3867 (
            .O(N__25375),
            .I(N__25369));
    Span12Mux_s3_h I__3866 (
            .O(N__25372),
            .I(N__25366));
    Sp12to4 I__3865 (
            .O(N__25369),
            .I(N__25361));
    Span12Mux_v I__3864 (
            .O(N__25366),
            .I(N__25361));
    Odrv12 I__3863 (
            .O(N__25361),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__3862 (
            .O(N__25358),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__3861 (
            .O(N__25355),
            .I(N__25351));
    InMux I__3860 (
            .O(N__25354),
            .I(N__25348));
    LocalMux I__3859 (
            .O(N__25351),
            .I(N__25345));
    LocalMux I__3858 (
            .O(N__25348),
            .I(N__25342));
    Span12Mux_s2_h I__3857 (
            .O(N__25345),
            .I(N__25339));
    Span4Mux_v I__3856 (
            .O(N__25342),
            .I(N__25336));
    Span12Mux_v I__3855 (
            .O(N__25339),
            .I(N__25333));
    Odrv4 I__3854 (
            .O(N__25336),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv12 I__3853 (
            .O(N__25333),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__3852 (
            .O(N__25328),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__3851 (
            .O(N__25325),
            .I(N__25321));
    InMux I__3850 (
            .O(N__25324),
            .I(N__25318));
    LocalMux I__3849 (
            .O(N__25321),
            .I(N__25315));
    LocalMux I__3848 (
            .O(N__25318),
            .I(N__25312));
    Span12Mux_s1_h I__3847 (
            .O(N__25315),
            .I(N__25309));
    Span4Mux_v I__3846 (
            .O(N__25312),
            .I(N__25306));
    Span12Mux_v I__3845 (
            .O(N__25309),
            .I(N__25303));
    Odrv4 I__3844 (
            .O(N__25306),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv12 I__3843 (
            .O(N__25303),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__3842 (
            .O(N__25298),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__3841 (
            .O(N__25295),
            .I(N__25291));
    InMux I__3840 (
            .O(N__25294),
            .I(N__25288));
    LocalMux I__3839 (
            .O(N__25291),
            .I(N__25285));
    LocalMux I__3838 (
            .O(N__25288),
            .I(N__25282));
    Span12Mux_s8_h I__3837 (
            .O(N__25285),
            .I(N__25279));
    Span4Mux_h I__3836 (
            .O(N__25282),
            .I(N__25276));
    Span12Mux_v I__3835 (
            .O(N__25279),
            .I(N__25273));
    Odrv4 I__3834 (
            .O(N__25276),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv12 I__3833 (
            .O(N__25273),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__3832 (
            .O(N__25268),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__3831 (
            .O(N__25265),
            .I(N__25262));
    LocalMux I__3830 (
            .O(N__25262),
            .I(N__25258));
    InMux I__3829 (
            .O(N__25261),
            .I(N__25255));
    Sp12to4 I__3828 (
            .O(N__25258),
            .I(N__25252));
    LocalMux I__3827 (
            .O(N__25255),
            .I(N__25249));
    Span12Mux_s11_h I__3826 (
            .O(N__25252),
            .I(N__25246));
    Span4Mux_h I__3825 (
            .O(N__25249),
            .I(N__25243));
    Span12Mux_v I__3824 (
            .O(N__25246),
            .I(N__25240));
    Odrv4 I__3823 (
            .O(N__25243),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv12 I__3822 (
            .O(N__25240),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__3821 (
            .O(N__25235),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__3820 (
            .O(N__25232),
            .I(N__25229));
    LocalMux I__3819 (
            .O(N__25229),
            .I(N__25225));
    InMux I__3818 (
            .O(N__25228),
            .I(N__25222));
    Sp12to4 I__3817 (
            .O(N__25225),
            .I(N__25219));
    LocalMux I__3816 (
            .O(N__25222),
            .I(N__25216));
    Span12Mux_s10_h I__3815 (
            .O(N__25219),
            .I(N__25213));
    Span4Mux_h I__3814 (
            .O(N__25216),
            .I(N__25210));
    Span12Mux_v I__3813 (
            .O(N__25213),
            .I(N__25207));
    Odrv4 I__3812 (
            .O(N__25210),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv12 I__3811 (
            .O(N__25207),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__3810 (
            .O(N__25202),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__3809 (
            .O(N__25199),
            .I(N__25196));
    LocalMux I__3808 (
            .O(N__25196),
            .I(N__25192));
    InMux I__3807 (
            .O(N__25195),
            .I(N__25189));
    Sp12to4 I__3806 (
            .O(N__25192),
            .I(N__25186));
    LocalMux I__3805 (
            .O(N__25189),
            .I(N__25183));
    Span12Mux_s5_h I__3804 (
            .O(N__25186),
            .I(N__25180));
    Span4Mux_h I__3803 (
            .O(N__25183),
            .I(N__25177));
    Span12Mux_v I__3802 (
            .O(N__25180),
            .I(N__25174));
    Odrv4 I__3801 (
            .O(N__25177),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv12 I__3800 (
            .O(N__25174),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__3799 (
            .O(N__25169),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__3798 (
            .O(N__25166),
            .I(N__25163));
    LocalMux I__3797 (
            .O(N__25163),
            .I(N__25160));
    Span4Mux_v I__3796 (
            .O(N__25160),
            .I(N__25156));
    InMux I__3795 (
            .O(N__25159),
            .I(N__25153));
    Sp12to4 I__3794 (
            .O(N__25156),
            .I(N__25150));
    LocalMux I__3793 (
            .O(N__25153),
            .I(N__25145));
    Span12Mux_s4_h I__3792 (
            .O(N__25150),
            .I(N__25145));
    Span12Mux_v I__3791 (
            .O(N__25145),
            .I(N__25142));
    Odrv12 I__3790 (
            .O(N__25142),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__3789 (
            .O(N__25139),
            .I(bfn_8_20_0_));
    InMux I__3788 (
            .O(N__25136),
            .I(N__25133));
    LocalMux I__3787 (
            .O(N__25133),
            .I(N__25129));
    InMux I__3786 (
            .O(N__25132),
            .I(N__25126));
    Span4Mux_v I__3785 (
            .O(N__25129),
            .I(N__25123));
    LocalMux I__3784 (
            .O(N__25126),
            .I(N__25120));
    Sp12to4 I__3783 (
            .O(N__25123),
            .I(N__25117));
    Span4Mux_h I__3782 (
            .O(N__25120),
            .I(N__25114));
    Span12Mux_s8_h I__3781 (
            .O(N__25117),
            .I(N__25111));
    Odrv4 I__3780 (
            .O(N__25114),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv12 I__3779 (
            .O(N__25111),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__3778 (
            .O(N__25106),
            .I(N__25100));
    InMux I__3777 (
            .O(N__25105),
            .I(N__25100));
    LocalMux I__3776 (
            .O(N__25100),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ));
    CascadeMux I__3775 (
            .O(N__25097),
            .I(N__25094));
    InMux I__3774 (
            .O(N__25094),
            .I(N__25087));
    InMux I__3773 (
            .O(N__25093),
            .I(N__25087));
    InMux I__3772 (
            .O(N__25092),
            .I(N__25084));
    LocalMux I__3771 (
            .O(N__25087),
            .I(N__25081));
    LocalMux I__3770 (
            .O(N__25084),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    Odrv12 I__3769 (
            .O(N__25081),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    CascadeMux I__3768 (
            .O(N__25076),
            .I(N__25072));
    InMux I__3767 (
            .O(N__25075),
            .I(N__25066));
    InMux I__3766 (
            .O(N__25072),
            .I(N__25066));
    InMux I__3765 (
            .O(N__25071),
            .I(N__25063));
    LocalMux I__3764 (
            .O(N__25066),
            .I(N__25060));
    LocalMux I__3763 (
            .O(N__25063),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    Odrv12 I__3762 (
            .O(N__25060),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    CascadeMux I__3761 (
            .O(N__25055),
            .I(N__25052));
    InMux I__3760 (
            .O(N__25052),
            .I(N__25049));
    LocalMux I__3759 (
            .O(N__25049),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt26 ));
    InMux I__3758 (
            .O(N__25046),
            .I(N__25043));
    LocalMux I__3757 (
            .O(N__25043),
            .I(N__25040));
    Span4Mux_h I__3756 (
            .O(N__25040),
            .I(N__25037));
    Odrv4 I__3755 (
            .O(N__25037),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    CascadeMux I__3754 (
            .O(N__25034),
            .I(N__25031));
    InMux I__3753 (
            .O(N__25031),
            .I(N__25025));
    InMux I__3752 (
            .O(N__25030),
            .I(N__25025));
    LocalMux I__3751 (
            .O(N__25025),
            .I(N__25022));
    Odrv4 I__3750 (
            .O(N__25022),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    CascadeMux I__3749 (
            .O(N__25019),
            .I(N__25016));
    InMux I__3748 (
            .O(N__25016),
            .I(N__25013));
    LocalMux I__3747 (
            .O(N__25013),
            .I(N__25009));
    InMux I__3746 (
            .O(N__25012),
            .I(N__25006));
    Span4Mux_h I__3745 (
            .O(N__25009),
            .I(N__25003));
    LocalMux I__3744 (
            .O(N__25006),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    Odrv4 I__3743 (
            .O(N__25003),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    InMux I__3742 (
            .O(N__24998),
            .I(N__24994));
    InMux I__3741 (
            .O(N__24997),
            .I(N__24991));
    LocalMux I__3740 (
            .O(N__24994),
            .I(N__24988));
    LocalMux I__3739 (
            .O(N__24991),
            .I(N__24985));
    Sp12to4 I__3738 (
            .O(N__24988),
            .I(N__24982));
    Span12Mux_v I__3737 (
            .O(N__24985),
            .I(N__24977));
    Span12Mux_v I__3736 (
            .O(N__24982),
            .I(N__24977));
    Odrv12 I__3735 (
            .O(N__24977),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__3734 (
            .O(N__24974),
            .I(N__24971));
    LocalMux I__3733 (
            .O(N__24971),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__3732 (
            .O(N__24968),
            .I(N__24965));
    LocalMux I__3731 (
            .O(N__24965),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt24 ));
    CascadeMux I__3730 (
            .O(N__24962),
            .I(N__24959));
    InMux I__3729 (
            .O(N__24959),
            .I(N__24956));
    LocalMux I__3728 (
            .O(N__24956),
            .I(N__24953));
    Odrv4 I__3727 (
            .O(N__24953),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ));
    InMux I__3726 (
            .O(N__24950),
            .I(N__24947));
    LocalMux I__3725 (
            .O(N__24947),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    CascadeMux I__3724 (
            .O(N__24944),
            .I(N__24941));
    InMux I__3723 (
            .O(N__24941),
            .I(N__24938));
    LocalMux I__3722 (
            .O(N__24938),
            .I(N__24934));
    InMux I__3721 (
            .O(N__24937),
            .I(N__24931));
    Odrv4 I__3720 (
            .O(N__24934),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    LocalMux I__3719 (
            .O(N__24931),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    InMux I__3718 (
            .O(N__24926),
            .I(N__24923));
    LocalMux I__3717 (
            .O(N__24923),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ));
    InMux I__3716 (
            .O(N__24920),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ));
    InMux I__3715 (
            .O(N__24917),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    InMux I__3714 (
            .O(N__24914),
            .I(N__24910));
    InMux I__3713 (
            .O(N__24913),
            .I(N__24907));
    LocalMux I__3712 (
            .O(N__24910),
            .I(N__24904));
    LocalMux I__3711 (
            .O(N__24907),
            .I(N__24901));
    Span4Mux_h I__3710 (
            .O(N__24904),
            .I(N__24898));
    Span4Mux_h I__3709 (
            .O(N__24901),
            .I(N__24895));
    Odrv4 I__3708 (
            .O(N__24898),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv4 I__3707 (
            .O(N__24895),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    CascadeMux I__3706 (
            .O(N__24890),
            .I(elapsed_time_ns_1_RNI58DN9_0_27_cascade_));
    InMux I__3705 (
            .O(N__24887),
            .I(N__24884));
    LocalMux I__3704 (
            .O(N__24884),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ));
    InMux I__3703 (
            .O(N__24881),
            .I(N__24877));
    InMux I__3702 (
            .O(N__24880),
            .I(N__24874));
    LocalMux I__3701 (
            .O(N__24877),
            .I(N__24871));
    LocalMux I__3700 (
            .O(N__24874),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv12 I__3699 (
            .O(N__24871),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__3698 (
            .O(N__24866),
            .I(N__24863));
    InMux I__3697 (
            .O(N__24863),
            .I(N__24860));
    LocalMux I__3696 (
            .O(N__24860),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__3695 (
            .O(N__24857),
            .I(N__24854));
    LocalMux I__3694 (
            .O(N__24854),
            .I(N__24850));
    InMux I__3693 (
            .O(N__24853),
            .I(N__24847));
    Span4Mux_v I__3692 (
            .O(N__24850),
            .I(N__24844));
    LocalMux I__3691 (
            .O(N__24847),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__3690 (
            .O(N__24844),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__3689 (
            .O(N__24839),
            .I(N__24836));
    InMux I__3688 (
            .O(N__24836),
            .I(N__24833));
    LocalMux I__3687 (
            .O(N__24833),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__3686 (
            .O(N__24830),
            .I(N__24826));
    InMux I__3685 (
            .O(N__24829),
            .I(N__24823));
    LocalMux I__3684 (
            .O(N__24826),
            .I(N__24820));
    LocalMux I__3683 (
            .O(N__24823),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv12 I__3682 (
            .O(N__24820),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__3681 (
            .O(N__24815),
            .I(N__24812));
    InMux I__3680 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__3679 (
            .O(N__24809),
            .I(N__24806));
    Odrv4 I__3678 (
            .O(N__24806),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__3677 (
            .O(N__24803),
            .I(N__24799));
    InMux I__3676 (
            .O(N__24802),
            .I(N__24796));
    LocalMux I__3675 (
            .O(N__24799),
            .I(N__24793));
    LocalMux I__3674 (
            .O(N__24796),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv12 I__3673 (
            .O(N__24793),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__3672 (
            .O(N__24788),
            .I(N__24785));
    LocalMux I__3671 (
            .O(N__24785),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__3670 (
            .O(N__24782),
            .I(N__24778));
    InMux I__3669 (
            .O(N__24781),
            .I(N__24775));
    LocalMux I__3668 (
            .O(N__24778),
            .I(N__24772));
    LocalMux I__3667 (
            .O(N__24775),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv12 I__3666 (
            .O(N__24772),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__3665 (
            .O(N__24767),
            .I(N__24764));
    InMux I__3664 (
            .O(N__24764),
            .I(N__24761));
    LocalMux I__3663 (
            .O(N__24761),
            .I(N__24758));
    Odrv4 I__3662 (
            .O(N__24758),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__3661 (
            .O(N__24755),
            .I(N__24752));
    LocalMux I__3660 (
            .O(N__24752),
            .I(N__24749));
    Span4Mux_v I__3659 (
            .O(N__24749),
            .I(N__24746));
    Odrv4 I__3658 (
            .O(N__24746),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    InMux I__3657 (
            .O(N__24743),
            .I(N__24740));
    LocalMux I__3656 (
            .O(N__24740),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ));
    CascadeMux I__3655 (
            .O(N__24737),
            .I(N__24734));
    InMux I__3654 (
            .O(N__24734),
            .I(N__24731));
    LocalMux I__3653 (
            .O(N__24731),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt20 ));
    InMux I__3652 (
            .O(N__24728),
            .I(N__24725));
    LocalMux I__3651 (
            .O(N__24725),
            .I(N__24721));
    InMux I__3650 (
            .O(N__24724),
            .I(N__24718));
    Span4Mux_v I__3649 (
            .O(N__24721),
            .I(N__24715));
    LocalMux I__3648 (
            .O(N__24718),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__3647 (
            .O(N__24715),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__3646 (
            .O(N__24710),
            .I(N__24707));
    InMux I__3645 (
            .O(N__24707),
            .I(N__24704));
    LocalMux I__3644 (
            .O(N__24704),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__3643 (
            .O(N__24701),
            .I(N__24697));
    InMux I__3642 (
            .O(N__24700),
            .I(N__24694));
    LocalMux I__3641 (
            .O(N__24697),
            .I(N__24691));
    LocalMux I__3640 (
            .O(N__24694),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv12 I__3639 (
            .O(N__24691),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__3638 (
            .O(N__24686),
            .I(N__24683));
    InMux I__3637 (
            .O(N__24683),
            .I(N__24680));
    LocalMux I__3636 (
            .O(N__24680),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    InMux I__3635 (
            .O(N__24677),
            .I(N__24674));
    LocalMux I__3634 (
            .O(N__24674),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__3633 (
            .O(N__24671),
            .I(N__24667));
    InMux I__3632 (
            .O(N__24670),
            .I(N__24664));
    LocalMux I__3631 (
            .O(N__24667),
            .I(N__24661));
    LocalMux I__3630 (
            .O(N__24664),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv12 I__3629 (
            .O(N__24661),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__3628 (
            .O(N__24656),
            .I(N__24653));
    LocalMux I__3627 (
            .O(N__24653),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__3626 (
            .O(N__24650),
            .I(N__24646));
    InMux I__3625 (
            .O(N__24649),
            .I(N__24643));
    LocalMux I__3624 (
            .O(N__24646),
            .I(N__24640));
    LocalMux I__3623 (
            .O(N__24643),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv12 I__3622 (
            .O(N__24640),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__3621 (
            .O(N__24635),
            .I(N__24632));
    InMux I__3620 (
            .O(N__24632),
            .I(N__24629));
    LocalMux I__3619 (
            .O(N__24629),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__3618 (
            .O(N__24626),
            .I(N__24622));
    InMux I__3617 (
            .O(N__24625),
            .I(N__24619));
    LocalMux I__3616 (
            .O(N__24622),
            .I(N__24616));
    LocalMux I__3615 (
            .O(N__24619),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv12 I__3614 (
            .O(N__24616),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__3613 (
            .O(N__24611),
            .I(N__24608));
    InMux I__3612 (
            .O(N__24608),
            .I(N__24605));
    LocalMux I__3611 (
            .O(N__24605),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    InMux I__3610 (
            .O(N__24602),
            .I(N__24598));
    InMux I__3609 (
            .O(N__24601),
            .I(N__24595));
    LocalMux I__3608 (
            .O(N__24598),
            .I(N__24592));
    LocalMux I__3607 (
            .O(N__24595),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv12 I__3606 (
            .O(N__24592),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    CascadeMux I__3605 (
            .O(N__24587),
            .I(N__24584));
    InMux I__3604 (
            .O(N__24584),
            .I(N__24581));
    LocalMux I__3603 (
            .O(N__24581),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__3602 (
            .O(N__24578),
            .I(N__24574));
    InMux I__3601 (
            .O(N__24577),
            .I(N__24571));
    LocalMux I__3600 (
            .O(N__24574),
            .I(N__24568));
    LocalMux I__3599 (
            .O(N__24571),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv12 I__3598 (
            .O(N__24568),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__3597 (
            .O(N__24563),
            .I(N__24560));
    InMux I__3596 (
            .O(N__24560),
            .I(N__24557));
    LocalMux I__3595 (
            .O(N__24557),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__3594 (
            .O(N__24554),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__3593 (
            .O(N__24551),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__3592 (
            .O(N__24548),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__3591 (
            .O(N__24545),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__3590 (
            .O(N__24542),
            .I(N__24532));
    InMux I__3589 (
            .O(N__24541),
            .I(N__24532));
    InMux I__3588 (
            .O(N__24540),
            .I(N__24532));
    InMux I__3587 (
            .O(N__24539),
            .I(N__24529));
    LocalMux I__3586 (
            .O(N__24532),
            .I(N__24526));
    LocalMux I__3585 (
            .O(N__24529),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    Odrv4 I__3584 (
            .O(N__24526),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    InMux I__3583 (
            .O(N__24521),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__3582 (
            .O(N__24518),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__3581 (
            .O(N__24515),
            .I(N__24505));
    InMux I__3580 (
            .O(N__24514),
            .I(N__24505));
    InMux I__3579 (
            .O(N__24513),
            .I(N__24505));
    InMux I__3578 (
            .O(N__24512),
            .I(N__24502));
    LocalMux I__3577 (
            .O(N__24505),
            .I(N__24499));
    LocalMux I__3576 (
            .O(N__24502),
            .I(N__24494));
    Span4Mux_v I__3575 (
            .O(N__24499),
            .I(N__24494));
    Odrv4 I__3574 (
            .O(N__24494),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    InMux I__3573 (
            .O(N__24491),
            .I(N__24488));
    LocalMux I__3572 (
            .O(N__24488),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__3571 (
            .O(N__24485),
            .I(N__24482));
    InMux I__3570 (
            .O(N__24482),
            .I(N__24479));
    LocalMux I__3569 (
            .O(N__24479),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__3568 (
            .O(N__24476),
            .I(N__24473));
    LocalMux I__3567 (
            .O(N__24473),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    InMux I__3566 (
            .O(N__24470),
            .I(N__24466));
    InMux I__3565 (
            .O(N__24469),
            .I(N__24463));
    LocalMux I__3564 (
            .O(N__24466),
            .I(N__24460));
    LocalMux I__3563 (
            .O(N__24463),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv12 I__3562 (
            .O(N__24460),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__3561 (
            .O(N__24455),
            .I(N__24452));
    InMux I__3560 (
            .O(N__24452),
            .I(N__24449));
    LocalMux I__3559 (
            .O(N__24449),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__3558 (
            .O(N__24446),
            .I(N__24443));
    LocalMux I__3557 (
            .O(N__24443),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__3556 (
            .O(N__24440),
            .I(N__24436));
    InMux I__3555 (
            .O(N__24439),
            .I(N__24433));
    LocalMux I__3554 (
            .O(N__24436),
            .I(N__24430));
    LocalMux I__3553 (
            .O(N__24433),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv12 I__3552 (
            .O(N__24430),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    CascadeMux I__3551 (
            .O(N__24425),
            .I(N__24422));
    InMux I__3550 (
            .O(N__24422),
            .I(N__24419));
    LocalMux I__3549 (
            .O(N__24419),
            .I(N__24416));
    Odrv4 I__3548 (
            .O(N__24416),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__3547 (
            .O(N__24413),
            .I(bfn_8_7_0_));
    InMux I__3546 (
            .O(N__24410),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__3545 (
            .O(N__24407),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__3544 (
            .O(N__24404),
            .I(N__24397));
    InMux I__3543 (
            .O(N__24403),
            .I(N__24397));
    InMux I__3542 (
            .O(N__24402),
            .I(N__24394));
    LocalMux I__3541 (
            .O(N__24397),
            .I(N__24391));
    LocalMux I__3540 (
            .O(N__24394),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__3539 (
            .O(N__24391),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__3538 (
            .O(N__24386),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    CascadeMux I__3537 (
            .O(N__24383),
            .I(N__24380));
    InMux I__3536 (
            .O(N__24380),
            .I(N__24374));
    InMux I__3535 (
            .O(N__24379),
            .I(N__24374));
    LocalMux I__3534 (
            .O(N__24374),
            .I(N__24370));
    InMux I__3533 (
            .O(N__24373),
            .I(N__24367));
    Span4Mux_h I__3532 (
            .O(N__24370),
            .I(N__24364));
    LocalMux I__3531 (
            .O(N__24367),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__3530 (
            .O(N__24364),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__3529 (
            .O(N__24359),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__3528 (
            .O(N__24356),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__3527 (
            .O(N__24353),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__3526 (
            .O(N__24350),
            .I(N__24347));
    LocalMux I__3525 (
            .O(N__24347),
            .I(N__24342));
    InMux I__3524 (
            .O(N__24346),
            .I(N__24339));
    InMux I__3523 (
            .O(N__24345),
            .I(N__24336));
    Span4Mux_v I__3522 (
            .O(N__24342),
            .I(N__24331));
    LocalMux I__3521 (
            .O(N__24339),
            .I(N__24331));
    LocalMux I__3520 (
            .O(N__24336),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__3519 (
            .O(N__24331),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__3518 (
            .O(N__24326),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    CascadeMux I__3517 (
            .O(N__24323),
            .I(N__24320));
    InMux I__3516 (
            .O(N__24320),
            .I(N__24317));
    LocalMux I__3515 (
            .O(N__24317),
            .I(N__24312));
    InMux I__3514 (
            .O(N__24316),
            .I(N__24309));
    InMux I__3513 (
            .O(N__24315),
            .I(N__24306));
    Span4Mux_v I__3512 (
            .O(N__24312),
            .I(N__24303));
    LocalMux I__3511 (
            .O(N__24309),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__3510 (
            .O(N__24306),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    Odrv4 I__3509 (
            .O(N__24303),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__3508 (
            .O(N__24296),
            .I(bfn_8_8_0_));
    InMux I__3507 (
            .O(N__24293),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__3506 (
            .O(N__24290),
            .I(bfn_8_6_0_));
    InMux I__3505 (
            .O(N__24287),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__3504 (
            .O(N__24284),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__3503 (
            .O(N__24281),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__3502 (
            .O(N__24278),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__3501 (
            .O(N__24275),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__3500 (
            .O(N__24272),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__3499 (
            .O(N__24269),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__3498 (
            .O(N__24266),
            .I(N__24263));
    LocalMux I__3497 (
            .O(N__24263),
            .I(N__24260));
    Odrv12 I__3496 (
            .O(N__24260),
            .I(il_max_comp1_c));
    InMux I__3495 (
            .O(N__24257),
            .I(N__24254));
    LocalMux I__3494 (
            .O(N__24254),
            .I(N__24251));
    Span4Mux_h I__3493 (
            .O(N__24251),
            .I(N__24248));
    Span4Mux_v I__3492 (
            .O(N__24248),
            .I(N__24245));
    Odrv4 I__3491 (
            .O(N__24245),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ));
    InMux I__3490 (
            .O(N__24242),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__3489 (
            .O(N__24239),
            .I(N__24236));
    InMux I__3488 (
            .O(N__24236),
            .I(N__24233));
    LocalMux I__3487 (
            .O(N__24233),
            .I(N__24230));
    Span4Mux_v I__3486 (
            .O(N__24230),
            .I(N__24227));
    Odrv4 I__3485 (
            .O(N__24227),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ));
    InMux I__3484 (
            .O(N__24224),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__3483 (
            .O(N__24221),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__3482 (
            .O(N__24218),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__3481 (
            .O(N__24215),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__3480 (
            .O(N__24212),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__3479 (
            .O(N__24209),
            .I(N__24206));
    LocalMux I__3478 (
            .O(N__24206),
            .I(N__24203));
    Span4Mux_h I__3477 (
            .O(N__24203),
            .I(N__24200));
    Odrv4 I__3476 (
            .O(N__24200),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__3475 (
            .O(N__24197),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__3474 (
            .O(N__24194),
            .I(N__24191));
    LocalMux I__3473 (
            .O(N__24191),
            .I(N__24188));
    Span4Mux_h I__3472 (
            .O(N__24188),
            .I(N__24185));
    Odrv4 I__3471 (
            .O(N__24185),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    InMux I__3470 (
            .O(N__24182),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    InMux I__3469 (
            .O(N__24179),
            .I(N__24176));
    LocalMux I__3468 (
            .O(N__24176),
            .I(N__24173));
    Span4Mux_v I__3467 (
            .O(N__24173),
            .I(N__24170));
    Odrv4 I__3466 (
            .O(N__24170),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    InMux I__3465 (
            .O(N__24167),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__3464 (
            .O(N__24164),
            .I(N__24161));
    LocalMux I__3463 (
            .O(N__24161),
            .I(N__24158));
    Span4Mux_h I__3462 (
            .O(N__24158),
            .I(N__24155));
    Odrv4 I__3461 (
            .O(N__24155),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__3460 (
            .O(N__24152),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__3459 (
            .O(N__24149),
            .I(N__24146));
    LocalMux I__3458 (
            .O(N__24146),
            .I(N__24143));
    Span4Mux_h I__3457 (
            .O(N__24143),
            .I(N__24140));
    Odrv4 I__3456 (
            .O(N__24140),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    InMux I__3455 (
            .O(N__24137),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    InMux I__3454 (
            .O(N__24134),
            .I(bfn_7_24_0_));
    InMux I__3453 (
            .O(N__24131),
            .I(N__24128));
    LocalMux I__3452 (
            .O(N__24128),
            .I(N__24125));
    Span4Mux_h I__3451 (
            .O(N__24125),
            .I(N__24122));
    Odrv4 I__3450 (
            .O(N__24122),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    InMux I__3449 (
            .O(N__24119),
            .I(N__24116));
    LocalMux I__3448 (
            .O(N__24116),
            .I(N__24113));
    Span4Mux_v I__3447 (
            .O(N__24113),
            .I(N__24110));
    Odrv4 I__3446 (
            .O(N__24110),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ));
    InMux I__3445 (
            .O(N__24107),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    InMux I__3444 (
            .O(N__24104),
            .I(N__24101));
    LocalMux I__3443 (
            .O(N__24101),
            .I(N__24096));
    InMux I__3442 (
            .O(N__24100),
            .I(N__24093));
    InMux I__3441 (
            .O(N__24099),
            .I(N__24090));
    Span4Mux_h I__3440 (
            .O(N__24096),
            .I(N__24087));
    LocalMux I__3439 (
            .O(N__24093),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__3438 (
            .O(N__24090),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    Odrv4 I__3437 (
            .O(N__24087),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    InMux I__3436 (
            .O(N__24080),
            .I(N__24076));
    InMux I__3435 (
            .O(N__24079),
            .I(N__24073));
    LocalMux I__3434 (
            .O(N__24076),
            .I(N__24070));
    LocalMux I__3433 (
            .O(N__24073),
            .I(N__24067));
    Span4Mux_h I__3432 (
            .O(N__24070),
            .I(N__24064));
    Span4Mux_v I__3431 (
            .O(N__24067),
            .I(N__24061));
    Odrv4 I__3430 (
            .O(N__24064),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    Odrv4 I__3429 (
            .O(N__24061),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    CascadeMux I__3428 (
            .O(N__24056),
            .I(N__24050));
    CascadeMux I__3427 (
            .O(N__24055),
            .I(N__24047));
    CascadeMux I__3426 (
            .O(N__24054),
            .I(N__24044));
    InMux I__3425 (
            .O(N__24053),
            .I(N__24041));
    InMux I__3424 (
            .O(N__24050),
            .I(N__24038));
    InMux I__3423 (
            .O(N__24047),
            .I(N__24035));
    InMux I__3422 (
            .O(N__24044),
            .I(N__24032));
    LocalMux I__3421 (
            .O(N__24041),
            .I(N__24027));
    LocalMux I__3420 (
            .O(N__24038),
            .I(N__24020));
    LocalMux I__3419 (
            .O(N__24035),
            .I(N__24020));
    LocalMux I__3418 (
            .O(N__24032),
            .I(N__24020));
    InMux I__3417 (
            .O(N__24031),
            .I(N__24015));
    CascadeMux I__3416 (
            .O(N__24030),
            .I(N__24012));
    Span4Mux_v I__3415 (
            .O(N__24027),
            .I(N__24004));
    Span4Mux_v I__3414 (
            .O(N__24020),
            .I(N__24004));
    InMux I__3413 (
            .O(N__24019),
            .I(N__24001));
    InMux I__3412 (
            .O(N__24018),
            .I(N__23998));
    LocalMux I__3411 (
            .O(N__24015),
            .I(N__23995));
    InMux I__3410 (
            .O(N__24012),
            .I(N__23986));
    InMux I__3409 (
            .O(N__24011),
            .I(N__23986));
    InMux I__3408 (
            .O(N__24010),
            .I(N__23986));
    InMux I__3407 (
            .O(N__24009),
            .I(N__23986));
    Odrv4 I__3406 (
            .O(N__24004),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    LocalMux I__3405 (
            .O(N__24001),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    LocalMux I__3404 (
            .O(N__23998),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__3403 (
            .O(N__23995),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    LocalMux I__3402 (
            .O(N__23986),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    InMux I__3401 (
            .O(N__23975),
            .I(N__23972));
    LocalMux I__3400 (
            .O(N__23972),
            .I(N__23969));
    Span4Mux_v I__3399 (
            .O(N__23969),
            .I(N__23966));
    Odrv4 I__3398 (
            .O(N__23966),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__3397 (
            .O(N__23963),
            .I(N__23960));
    LocalMux I__3396 (
            .O(N__23960),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__3395 (
            .O(N__23957),
            .I(N__23954));
    LocalMux I__3394 (
            .O(N__23954),
            .I(N__23950));
    InMux I__3393 (
            .O(N__23953),
            .I(N__23947));
    Odrv12 I__3392 (
            .O(N__23950),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    LocalMux I__3391 (
            .O(N__23947),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    CascadeMux I__3390 (
            .O(N__23942),
            .I(N__23937));
    CascadeMux I__3389 (
            .O(N__23941),
            .I(N__23934));
    CascadeMux I__3388 (
            .O(N__23940),
            .I(N__23931));
    InMux I__3387 (
            .O(N__23937),
            .I(N__23924));
    InMux I__3386 (
            .O(N__23934),
            .I(N__23924));
    InMux I__3385 (
            .O(N__23931),
            .I(N__23924));
    LocalMux I__3384 (
            .O(N__23924),
            .I(N__23921));
    Odrv4 I__3383 (
            .O(N__23921),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    InMux I__3382 (
            .O(N__23918),
            .I(N__23912));
    InMux I__3381 (
            .O(N__23917),
            .I(N__23909));
    InMux I__3380 (
            .O(N__23916),
            .I(N__23904));
    InMux I__3379 (
            .O(N__23915),
            .I(N__23904));
    LocalMux I__3378 (
            .O(N__23912),
            .I(N__23896));
    LocalMux I__3377 (
            .O(N__23909),
            .I(N__23896));
    LocalMux I__3376 (
            .O(N__23904),
            .I(N__23896));
    InMux I__3375 (
            .O(N__23903),
            .I(N__23893));
    Span4Mux_v I__3374 (
            .O(N__23896),
            .I(N__23890));
    LocalMux I__3373 (
            .O(N__23893),
            .I(N__23887));
    Span4Mux_v I__3372 (
            .O(N__23890),
            .I(N__23884));
    Odrv12 I__3371 (
            .O(N__23887),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__3370 (
            .O(N__23884),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__3369 (
            .O(N__23879),
            .I(N__23876));
    LocalMux I__3368 (
            .O(N__23876),
            .I(N__23873));
    Span4Mux_h I__3367 (
            .O(N__23873),
            .I(N__23870));
    Odrv4 I__3366 (
            .O(N__23870),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    InMux I__3365 (
            .O(N__23867),
            .I(N__23864));
    LocalMux I__3364 (
            .O(N__23864),
            .I(N__23861));
    Span4Mux_h I__3363 (
            .O(N__23861),
            .I(N__23858));
    Odrv4 I__3362 (
            .O(N__23858),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__3361 (
            .O(N__23855),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    InMux I__3360 (
            .O(N__23852),
            .I(N__23849));
    LocalMux I__3359 (
            .O(N__23849),
            .I(N__23846));
    Span4Mux_h I__3358 (
            .O(N__23846),
            .I(N__23843));
    Odrv4 I__3357 (
            .O(N__23843),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    InMux I__3356 (
            .O(N__23840),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__3355 (
            .O(N__23837),
            .I(N__23831));
    InMux I__3354 (
            .O(N__23836),
            .I(N__23831));
    LocalMux I__3353 (
            .O(N__23831),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    CascadeMux I__3352 (
            .O(N__23828),
            .I(\phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ));
    CascadeMux I__3351 (
            .O(N__23825),
            .I(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ));
    CascadeMux I__3350 (
            .O(N__23822),
            .I(elapsed_time_ns_1_RNIH33T9_0_5_cascade_));
    InMux I__3349 (
            .O(N__23819),
            .I(N__23814));
    InMux I__3348 (
            .O(N__23818),
            .I(N__23811));
    InMux I__3347 (
            .O(N__23817),
            .I(N__23808));
    LocalMux I__3346 (
            .O(N__23814),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    LocalMux I__3345 (
            .O(N__23811),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    LocalMux I__3344 (
            .O(N__23808),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    InMux I__3343 (
            .O(N__23801),
            .I(N__23798));
    LocalMux I__3342 (
            .O(N__23798),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    InMux I__3341 (
            .O(N__23795),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    CascadeMux I__3340 (
            .O(N__23792),
            .I(N__23787));
    InMux I__3339 (
            .O(N__23791),
            .I(N__23784));
    InMux I__3338 (
            .O(N__23790),
            .I(N__23781));
    InMux I__3337 (
            .O(N__23787),
            .I(N__23778));
    LocalMux I__3336 (
            .O(N__23784),
            .I(N__23775));
    LocalMux I__3335 (
            .O(N__23781),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    LocalMux I__3334 (
            .O(N__23778),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__3333 (
            .O(N__23775),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__3332 (
            .O(N__23768),
            .I(N__23765));
    LocalMux I__3331 (
            .O(N__23765),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    InMux I__3330 (
            .O(N__23762),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    InMux I__3329 (
            .O(N__23759),
            .I(N__23754));
    InMux I__3328 (
            .O(N__23758),
            .I(N__23751));
    InMux I__3327 (
            .O(N__23757),
            .I(N__23748));
    LocalMux I__3326 (
            .O(N__23754),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__3325 (
            .O(N__23751),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__3324 (
            .O(N__23748),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    InMux I__3323 (
            .O(N__23741),
            .I(N__23738));
    LocalMux I__3322 (
            .O(N__23738),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    InMux I__3321 (
            .O(N__23735),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    InMux I__3320 (
            .O(N__23732),
            .I(N__23728));
    InMux I__3319 (
            .O(N__23731),
            .I(N__23725));
    LocalMux I__3318 (
            .O(N__23728),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__3317 (
            .O(N__23725),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    InMux I__3316 (
            .O(N__23720),
            .I(N__23717));
    LocalMux I__3315 (
            .O(N__23717),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__3314 (
            .O(N__23714),
            .I(bfn_5_27_0_));
    InMux I__3313 (
            .O(N__23711),
            .I(N__23706));
    InMux I__3312 (
            .O(N__23710),
            .I(N__23703));
    InMux I__3311 (
            .O(N__23709),
            .I(N__23700));
    LocalMux I__3310 (
            .O(N__23706),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    LocalMux I__3309 (
            .O(N__23703),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    LocalMux I__3308 (
            .O(N__23700),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__3307 (
            .O(N__23693),
            .I(N__23690));
    LocalMux I__3306 (
            .O(N__23690),
            .I(N__23687));
    Odrv4 I__3305 (
            .O(N__23687),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__3304 (
            .O(N__23684),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__3303 (
            .O(N__23681),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__3302 (
            .O(N__23678),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__3301 (
            .O(N__23675),
            .I(N__23672));
    LocalMux I__3300 (
            .O(N__23672),
            .I(N__23669));
    Span4Mux_h I__3299 (
            .O(N__23669),
            .I(N__23666));
    Span4Mux_h I__3298 (
            .O(N__23666),
            .I(N__23663));
    Odrv4 I__3297 (
            .O(N__23663),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__3296 (
            .O(N__23660),
            .I(N__23657));
    LocalMux I__3295 (
            .O(N__23657),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__3294 (
            .O(N__23654),
            .I(N__23651));
    LocalMux I__3293 (
            .O(N__23651),
            .I(N__23648));
    Span4Mux_h I__3292 (
            .O(N__23648),
            .I(N__23645));
    Span4Mux_h I__3291 (
            .O(N__23645),
            .I(N__23642));
    Odrv4 I__3290 (
            .O(N__23642),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__3289 (
            .O(N__23639),
            .I(N__23636));
    LocalMux I__3288 (
            .O(N__23636),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    InMux I__3287 (
            .O(N__23633),
            .I(N__23630));
    LocalMux I__3286 (
            .O(N__23630),
            .I(N__23627));
    Span4Mux_v I__3285 (
            .O(N__23627),
            .I(N__23624));
    Span4Mux_h I__3284 (
            .O(N__23624),
            .I(N__23621));
    Odrv4 I__3283 (
            .O(N__23621),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__3282 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__3281 (
            .O(N__23615),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__3280 (
            .O(N__23612),
            .I(N__23609));
    LocalMux I__3279 (
            .O(N__23609),
            .I(N__23606));
    Span4Mux_h I__3278 (
            .O(N__23606),
            .I(N__23603));
    Span4Mux_h I__3277 (
            .O(N__23603),
            .I(N__23600));
    Odrv4 I__3276 (
            .O(N__23600),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__3275 (
            .O(N__23597),
            .I(N__23594));
    LocalMux I__3274 (
            .O(N__23594),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__3273 (
            .O(N__23591),
            .I(N__23588));
    LocalMux I__3272 (
            .O(N__23588),
            .I(N__23585));
    Span4Mux_h I__3271 (
            .O(N__23585),
            .I(N__23582));
    Span4Mux_h I__3270 (
            .O(N__23582),
            .I(N__23579));
    Odrv4 I__3269 (
            .O(N__23579),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__3268 (
            .O(N__23576),
            .I(N__23573));
    LocalMux I__3267 (
            .O(N__23573),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__3266 (
            .O(N__23570),
            .I(N__23566));
    InMux I__3265 (
            .O(N__23569),
            .I(N__23562));
    LocalMux I__3264 (
            .O(N__23566),
            .I(N__23559));
    InMux I__3263 (
            .O(N__23565),
            .I(N__23556));
    LocalMux I__3262 (
            .O(N__23562),
            .I(N__23553));
    Span4Mux_h I__3261 (
            .O(N__23559),
            .I(N__23550));
    LocalMux I__3260 (
            .O(N__23556),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__3259 (
            .O(N__23553),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__3258 (
            .O(N__23550),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    InMux I__3257 (
            .O(N__23543),
            .I(N__23540));
    LocalMux I__3256 (
            .O(N__23540),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    InMux I__3255 (
            .O(N__23537),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    InMux I__3254 (
            .O(N__23534),
            .I(N__23531));
    LocalMux I__3253 (
            .O(N__23531),
            .I(N__23527));
    InMux I__3252 (
            .O(N__23530),
            .I(N__23524));
    Span12Mux_s6_v I__3251 (
            .O(N__23527),
            .I(N__23521));
    LocalMux I__3250 (
            .O(N__23524),
            .I(N__23518));
    Odrv12 I__3249 (
            .O(N__23521),
            .I(\pwm_generator_inst.un3_threshold ));
    Odrv4 I__3248 (
            .O(N__23518),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__3247 (
            .O(N__23513),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    InMux I__3246 (
            .O(N__23510),
            .I(N__23506));
    InMux I__3245 (
            .O(N__23509),
            .I(N__23502));
    LocalMux I__3244 (
            .O(N__23506),
            .I(N__23499));
    InMux I__3243 (
            .O(N__23505),
            .I(N__23496));
    LocalMux I__3242 (
            .O(N__23502),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv4 I__3241 (
            .O(N__23499),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__3240 (
            .O(N__23496),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__3239 (
            .O(N__23489),
            .I(N__23486));
    LocalMux I__3238 (
            .O(N__23486),
            .I(N__23483));
    Odrv4 I__3237 (
            .O(N__23483),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    InMux I__3236 (
            .O(N__23480),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__3235 (
            .O(N__23477),
            .I(N__23474));
    LocalMux I__3234 (
            .O(N__23474),
            .I(N__23471));
    Span4Mux_h I__3233 (
            .O(N__23471),
            .I(N__23468));
    Sp12to4 I__3232 (
            .O(N__23468),
            .I(N__23465));
    Span12Mux_s5_v I__3231 (
            .O(N__23465),
            .I(N__23462));
    Span12Mux_h I__3230 (
            .O(N__23462),
            .I(N__23459));
    Odrv12 I__3229 (
            .O(N__23459),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__3228 (
            .O(N__23456),
            .I(N__23453));
    LocalMux I__3227 (
            .O(N__23453),
            .I(N__23450));
    Span4Mux_h I__3226 (
            .O(N__23450),
            .I(N__23447));
    Odrv4 I__3225 (
            .O(N__23447),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    CascadeMux I__3224 (
            .O(N__23444),
            .I(N__23440));
    InMux I__3223 (
            .O(N__23443),
            .I(N__23437));
    InMux I__3222 (
            .O(N__23440),
            .I(N__23434));
    LocalMux I__3221 (
            .O(N__23437),
            .I(N__23431));
    LocalMux I__3220 (
            .O(N__23434),
            .I(N__23428));
    Span4Mux_h I__3219 (
            .O(N__23431),
            .I(N__23425));
    Odrv4 I__3218 (
            .O(N__23428),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    Odrv4 I__3217 (
            .O(N__23425),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    InMux I__3216 (
            .O(N__23420),
            .I(N__23416));
    InMux I__3215 (
            .O(N__23419),
            .I(N__23413));
    LocalMux I__3214 (
            .O(N__23416),
            .I(N__23410));
    LocalMux I__3213 (
            .O(N__23413),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    Odrv4 I__3212 (
            .O(N__23410),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    InMux I__3211 (
            .O(N__23405),
            .I(N__23402));
    LocalMux I__3210 (
            .O(N__23402),
            .I(N__23399));
    Span4Mux_h I__3209 (
            .O(N__23399),
            .I(N__23396));
    Span4Mux_h I__3208 (
            .O(N__23396),
            .I(N__23393));
    Odrv4 I__3207 (
            .O(N__23393),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__3206 (
            .O(N__23390),
            .I(N__23387));
    LocalMux I__3205 (
            .O(N__23387),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__3204 (
            .O(N__23384),
            .I(N__23381));
    LocalMux I__3203 (
            .O(N__23381),
            .I(N__23378));
    Span4Mux_h I__3202 (
            .O(N__23378),
            .I(N__23375));
    Span4Mux_h I__3201 (
            .O(N__23375),
            .I(N__23372));
    Odrv4 I__3200 (
            .O(N__23372),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__3199 (
            .O(N__23369),
            .I(N__23366));
    LocalMux I__3198 (
            .O(N__23366),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__3197 (
            .O(N__23363),
            .I(N__23360));
    LocalMux I__3196 (
            .O(N__23360),
            .I(N__23357));
    Span12Mux_h I__3195 (
            .O(N__23357),
            .I(N__23354));
    Odrv12 I__3194 (
            .O(N__23354),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__3193 (
            .O(N__23351),
            .I(N__23348));
    LocalMux I__3192 (
            .O(N__23348),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__3191 (
            .O(N__23345),
            .I(N__23342));
    LocalMux I__3190 (
            .O(N__23342),
            .I(N__23339));
    Span12Mux_s7_v I__3189 (
            .O(N__23339),
            .I(N__23336));
    Odrv12 I__3188 (
            .O(N__23336),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__3187 (
            .O(N__23333),
            .I(N__23330));
    LocalMux I__3186 (
            .O(N__23330),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__3185 (
            .O(N__23327),
            .I(N__23324));
    LocalMux I__3184 (
            .O(N__23324),
            .I(N__23321));
    Span4Mux_h I__3183 (
            .O(N__23321),
            .I(N__23318));
    Span4Mux_h I__3182 (
            .O(N__23318),
            .I(N__23315));
    Odrv4 I__3181 (
            .O(N__23315),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__3180 (
            .O(N__23312),
            .I(N__23309));
    LocalMux I__3179 (
            .O(N__23309),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    CascadeMux I__3178 (
            .O(N__23306),
            .I(N__23303));
    InMux I__3177 (
            .O(N__23303),
            .I(N__23300));
    LocalMux I__3176 (
            .O(N__23300),
            .I(N__23297));
    Odrv4 I__3175 (
            .O(N__23297),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    CascadeMux I__3174 (
            .O(N__23294),
            .I(N__23291));
    InMux I__3173 (
            .O(N__23291),
            .I(N__23288));
    LocalMux I__3172 (
            .O(N__23288),
            .I(N__23284));
    InMux I__3171 (
            .O(N__23287),
            .I(N__23279));
    Span4Mux_v I__3170 (
            .O(N__23284),
            .I(N__23276));
    InMux I__3169 (
            .O(N__23283),
            .I(N__23271));
    InMux I__3168 (
            .O(N__23282),
            .I(N__23271));
    LocalMux I__3167 (
            .O(N__23279),
            .I(N__23268));
    Odrv4 I__3166 (
            .O(N__23276),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__3165 (
            .O(N__23271),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__3164 (
            .O(N__23268),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__3163 (
            .O(N__23261),
            .I(N__23249));
    InMux I__3162 (
            .O(N__23260),
            .I(N__23246));
    CascadeMux I__3161 (
            .O(N__23259),
            .I(N__23242));
    CascadeMux I__3160 (
            .O(N__23258),
            .I(N__23239));
    CascadeMux I__3159 (
            .O(N__23257),
            .I(N__23236));
    InMux I__3158 (
            .O(N__23256),
            .I(N__23224));
    InMux I__3157 (
            .O(N__23255),
            .I(N__23217));
    InMux I__3156 (
            .O(N__23254),
            .I(N__23217));
    InMux I__3155 (
            .O(N__23253),
            .I(N__23212));
    InMux I__3154 (
            .O(N__23252),
            .I(N__23212));
    LocalMux I__3153 (
            .O(N__23249),
            .I(N__23207));
    LocalMux I__3152 (
            .O(N__23246),
            .I(N__23207));
    InMux I__3151 (
            .O(N__23245),
            .I(N__23204));
    InMux I__3150 (
            .O(N__23242),
            .I(N__23193));
    InMux I__3149 (
            .O(N__23239),
            .I(N__23193));
    InMux I__3148 (
            .O(N__23236),
            .I(N__23193));
    InMux I__3147 (
            .O(N__23235),
            .I(N__23193));
    InMux I__3146 (
            .O(N__23234),
            .I(N__23193));
    InMux I__3145 (
            .O(N__23233),
            .I(N__23190));
    InMux I__3144 (
            .O(N__23232),
            .I(N__23168));
    InMux I__3143 (
            .O(N__23231),
            .I(N__23168));
    InMux I__3142 (
            .O(N__23230),
            .I(N__23168));
    InMux I__3141 (
            .O(N__23229),
            .I(N__23168));
    InMux I__3140 (
            .O(N__23228),
            .I(N__23168));
    InMux I__3139 (
            .O(N__23227),
            .I(N__23168));
    LocalMux I__3138 (
            .O(N__23224),
            .I(N__23165));
    InMux I__3137 (
            .O(N__23223),
            .I(N__23160));
    InMux I__3136 (
            .O(N__23222),
            .I(N__23160));
    LocalMux I__3135 (
            .O(N__23217),
            .I(N__23156));
    LocalMux I__3134 (
            .O(N__23212),
            .I(N__23149));
    Span4Mux_h I__3133 (
            .O(N__23207),
            .I(N__23149));
    LocalMux I__3132 (
            .O(N__23204),
            .I(N__23149));
    LocalMux I__3131 (
            .O(N__23193),
            .I(N__23144));
    LocalMux I__3130 (
            .O(N__23190),
            .I(N__23144));
    InMux I__3129 (
            .O(N__23189),
            .I(N__23141));
    InMux I__3128 (
            .O(N__23188),
            .I(N__23128));
    InMux I__3127 (
            .O(N__23187),
            .I(N__23128));
    InMux I__3126 (
            .O(N__23186),
            .I(N__23128));
    InMux I__3125 (
            .O(N__23185),
            .I(N__23128));
    InMux I__3124 (
            .O(N__23184),
            .I(N__23128));
    InMux I__3123 (
            .O(N__23183),
            .I(N__23128));
    InMux I__3122 (
            .O(N__23182),
            .I(N__23123));
    InMux I__3121 (
            .O(N__23181),
            .I(N__23123));
    LocalMux I__3120 (
            .O(N__23168),
            .I(N__23120));
    Span4Mux_v I__3119 (
            .O(N__23165),
            .I(N__23117));
    LocalMux I__3118 (
            .O(N__23160),
            .I(N__23114));
    InMux I__3117 (
            .O(N__23159),
            .I(N__23111));
    Span4Mux_v I__3116 (
            .O(N__23156),
            .I(N__23106));
    Span4Mux_v I__3115 (
            .O(N__23149),
            .I(N__23106));
    Span4Mux_h I__3114 (
            .O(N__23144),
            .I(N__23103));
    LocalMux I__3113 (
            .O(N__23141),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3112 (
            .O(N__23128),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3111 (
            .O(N__23123),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3110 (
            .O(N__23120),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3109 (
            .O(N__23117),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv12 I__3108 (
            .O(N__23114),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__3107 (
            .O(N__23111),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3106 (
            .O(N__23106),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__3105 (
            .O(N__23103),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    CascadeMux I__3104 (
            .O(N__23084),
            .I(N__23078));
    InMux I__3103 (
            .O(N__23083),
            .I(N__23068));
    InMux I__3102 (
            .O(N__23082),
            .I(N__23068));
    InMux I__3101 (
            .O(N__23081),
            .I(N__23065));
    InMux I__3100 (
            .O(N__23078),
            .I(N__23058));
    InMux I__3099 (
            .O(N__23077),
            .I(N__23058));
    InMux I__3098 (
            .O(N__23076),
            .I(N__23055));
    InMux I__3097 (
            .O(N__23075),
            .I(N__23030));
    InMux I__3096 (
            .O(N__23074),
            .I(N__23030));
    InMux I__3095 (
            .O(N__23073),
            .I(N__23027));
    LocalMux I__3094 (
            .O(N__23068),
            .I(N__23024));
    LocalMux I__3093 (
            .O(N__23065),
            .I(N__23021));
    InMux I__3092 (
            .O(N__23064),
            .I(N__23016));
    InMux I__3091 (
            .O(N__23063),
            .I(N__23016));
    LocalMux I__3090 (
            .O(N__23058),
            .I(N__23011));
    LocalMux I__3089 (
            .O(N__23055),
            .I(N__23011));
    InMux I__3088 (
            .O(N__23054),
            .I(N__23002));
    InMux I__3087 (
            .O(N__23053),
            .I(N__23002));
    InMux I__3086 (
            .O(N__23052),
            .I(N__23002));
    InMux I__3085 (
            .O(N__23051),
            .I(N__23002));
    InMux I__3084 (
            .O(N__23050),
            .I(N__22997));
    InMux I__3083 (
            .O(N__23049),
            .I(N__22997));
    InMux I__3082 (
            .O(N__23048),
            .I(N__22990));
    InMux I__3081 (
            .O(N__23047),
            .I(N__22990));
    InMux I__3080 (
            .O(N__23046),
            .I(N__22990));
    InMux I__3079 (
            .O(N__23045),
            .I(N__22977));
    InMux I__3078 (
            .O(N__23044),
            .I(N__22977));
    InMux I__3077 (
            .O(N__23043),
            .I(N__22977));
    InMux I__3076 (
            .O(N__23042),
            .I(N__22977));
    InMux I__3075 (
            .O(N__23041),
            .I(N__22977));
    InMux I__3074 (
            .O(N__23040),
            .I(N__22977));
    InMux I__3073 (
            .O(N__23039),
            .I(N__22966));
    InMux I__3072 (
            .O(N__23038),
            .I(N__22966));
    InMux I__3071 (
            .O(N__23037),
            .I(N__22966));
    InMux I__3070 (
            .O(N__23036),
            .I(N__22966));
    InMux I__3069 (
            .O(N__23035),
            .I(N__22966));
    LocalMux I__3068 (
            .O(N__23030),
            .I(N__22963));
    LocalMux I__3067 (
            .O(N__23027),
            .I(N__22960));
    Span4Mux_v I__3066 (
            .O(N__23024),
            .I(N__22955));
    Span4Mux_v I__3065 (
            .O(N__23021),
            .I(N__22955));
    LocalMux I__3064 (
            .O(N__23016),
            .I(N__22950));
    Span4Mux_v I__3063 (
            .O(N__23011),
            .I(N__22950));
    LocalMux I__3062 (
            .O(N__23002),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    LocalMux I__3061 (
            .O(N__22997),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    LocalMux I__3060 (
            .O(N__22990),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    LocalMux I__3059 (
            .O(N__22977),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    LocalMux I__3058 (
            .O(N__22966),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__3057 (
            .O(N__22963),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv12 I__3056 (
            .O(N__22960),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__3055 (
            .O(N__22955),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    Odrv4 I__3054 (
            .O(N__22950),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    CascadeMux I__3053 (
            .O(N__22931),
            .I(N__22928));
    InMux I__3052 (
            .O(N__22928),
            .I(N__22925));
    LocalMux I__3051 (
            .O(N__22925),
            .I(N__22922));
    Span4Mux_h I__3050 (
            .O(N__22922),
            .I(N__22919));
    Odrv4 I__3049 (
            .O(N__22919),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    CascadeMux I__3048 (
            .O(N__22916),
            .I(N__22913));
    InMux I__3047 (
            .O(N__22913),
            .I(N__22909));
    InMux I__3046 (
            .O(N__22912),
            .I(N__22905));
    LocalMux I__3045 (
            .O(N__22909),
            .I(N__22901));
    CascadeMux I__3044 (
            .O(N__22908),
            .I(N__22898));
    LocalMux I__3043 (
            .O(N__22905),
            .I(N__22895));
    InMux I__3042 (
            .O(N__22904),
            .I(N__22892));
    Span4Mux_h I__3041 (
            .O(N__22901),
            .I(N__22889));
    InMux I__3040 (
            .O(N__22898),
            .I(N__22886));
    Span4Mux_h I__3039 (
            .O(N__22895),
            .I(N__22883));
    LocalMux I__3038 (
            .O(N__22892),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__3037 (
            .O(N__22889),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__3036 (
            .O(N__22886),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__3035 (
            .O(N__22883),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    CascadeMux I__3034 (
            .O(N__22874),
            .I(N__22870));
    InMux I__3033 (
            .O(N__22873),
            .I(N__22866));
    InMux I__3032 (
            .O(N__22870),
            .I(N__22863));
    InMux I__3031 (
            .O(N__22869),
            .I(N__22859));
    LocalMux I__3030 (
            .O(N__22866),
            .I(N__22854));
    LocalMux I__3029 (
            .O(N__22863),
            .I(N__22854));
    InMux I__3028 (
            .O(N__22862),
            .I(N__22851));
    LocalMux I__3027 (
            .O(N__22859),
            .I(N__22848));
    Span4Mux_v I__3026 (
            .O(N__22854),
            .I(N__22843));
    LocalMux I__3025 (
            .O(N__22851),
            .I(N__22843));
    Span4Mux_v I__3024 (
            .O(N__22848),
            .I(N__22840));
    Span4Mux_h I__3023 (
            .O(N__22843),
            .I(N__22837));
    Odrv4 I__3022 (
            .O(N__22840),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv4 I__3021 (
            .O(N__22837),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    InMux I__3020 (
            .O(N__22832),
            .I(N__22827));
    InMux I__3019 (
            .O(N__22831),
            .I(N__22824));
    InMux I__3018 (
            .O(N__22830),
            .I(N__22821));
    LocalMux I__3017 (
            .O(N__22827),
            .I(N__22817));
    LocalMux I__3016 (
            .O(N__22824),
            .I(N__22814));
    LocalMux I__3015 (
            .O(N__22821),
            .I(N__22811));
    InMux I__3014 (
            .O(N__22820),
            .I(N__22808));
    Span4Mux_h I__3013 (
            .O(N__22817),
            .I(N__22805));
    Span4Mux_v I__3012 (
            .O(N__22814),
            .I(N__22800));
    Span4Mux_h I__3011 (
            .O(N__22811),
            .I(N__22800));
    LocalMux I__3010 (
            .O(N__22808),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__3009 (
            .O(N__22805),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__3008 (
            .O(N__22800),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    CascadeMux I__3007 (
            .O(N__22793),
            .I(N__22788));
    CascadeMux I__3006 (
            .O(N__22792),
            .I(N__22785));
    InMux I__3005 (
            .O(N__22791),
            .I(N__22782));
    InMux I__3004 (
            .O(N__22788),
            .I(N__22779));
    InMux I__3003 (
            .O(N__22785),
            .I(N__22776));
    LocalMux I__3002 (
            .O(N__22782),
            .I(N__22773));
    LocalMux I__3001 (
            .O(N__22779),
            .I(N__22770));
    LocalMux I__3000 (
            .O(N__22776),
            .I(N__22767));
    Span4Mux_h I__2999 (
            .O(N__22773),
            .I(N__22763));
    Span4Mux_h I__2998 (
            .O(N__22770),
            .I(N__22758));
    Span4Mux_v I__2997 (
            .O(N__22767),
            .I(N__22758));
    InMux I__2996 (
            .O(N__22766),
            .I(N__22755));
    Odrv4 I__2995 (
            .O(N__22763),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__2994 (
            .O(N__22758),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__2993 (
            .O(N__22755),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__2992 (
            .O(N__22748),
            .I(N__22745));
    LocalMux I__2991 (
            .O(N__22745),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ));
    CascadeMux I__2990 (
            .O(N__22742),
            .I(N__22739));
    InMux I__2989 (
            .O(N__22739),
            .I(N__22736));
    LocalMux I__2988 (
            .O(N__22736),
            .I(N__22733));
    Span4Mux_h I__2987 (
            .O(N__22733),
            .I(N__22728));
    InMux I__2986 (
            .O(N__22732),
            .I(N__22724));
    InMux I__2985 (
            .O(N__22731),
            .I(N__22721));
    Span4Mux_v I__2984 (
            .O(N__22728),
            .I(N__22718));
    InMux I__2983 (
            .O(N__22727),
            .I(N__22715));
    LocalMux I__2982 (
            .O(N__22724),
            .I(N__22710));
    LocalMux I__2981 (
            .O(N__22721),
            .I(N__22710));
    Odrv4 I__2980 (
            .O(N__22718),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    LocalMux I__2979 (
            .O(N__22715),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv12 I__2978 (
            .O(N__22710),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__2977 (
            .O(N__22703),
            .I(N__22700));
    InMux I__2976 (
            .O(N__22700),
            .I(N__22696));
    InMux I__2975 (
            .O(N__22699),
            .I(N__22691));
    LocalMux I__2974 (
            .O(N__22696),
            .I(N__22688));
    InMux I__2973 (
            .O(N__22695),
            .I(N__22685));
    InMux I__2972 (
            .O(N__22694),
            .I(N__22682));
    LocalMux I__2971 (
            .O(N__22691),
            .I(N__22679));
    Odrv12 I__2970 (
            .O(N__22688),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__2969 (
            .O(N__22685),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__2968 (
            .O(N__22682),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__2967 (
            .O(N__22679),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    CascadeMux I__2966 (
            .O(N__22670),
            .I(\current_shift_inst.PI_CTRL.N_44_cascade_ ));
    InMux I__2965 (
            .O(N__22667),
            .I(N__22664));
    LocalMux I__2964 (
            .O(N__22664),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    InMux I__2963 (
            .O(N__22661),
            .I(N__22658));
    LocalMux I__2962 (
            .O(N__22658),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    InMux I__2961 (
            .O(N__22655),
            .I(N__22652));
    LocalMux I__2960 (
            .O(N__22652),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ));
    CascadeMux I__2959 (
            .O(N__22649),
            .I(N__22646));
    InMux I__2958 (
            .O(N__22646),
            .I(N__22643));
    LocalMux I__2957 (
            .O(N__22643),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    InMux I__2956 (
            .O(N__22640),
            .I(N__22637));
    LocalMux I__2955 (
            .O(N__22637),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    CascadeMux I__2954 (
            .O(N__22634),
            .I(N__22621));
    CascadeMux I__2953 (
            .O(N__22633),
            .I(N__22618));
    CascadeMux I__2952 (
            .O(N__22632),
            .I(N__22603));
    CascadeMux I__2951 (
            .O(N__22631),
            .I(N__22599));
    InMux I__2950 (
            .O(N__22630),
            .I(N__22582));
    InMux I__2949 (
            .O(N__22629),
            .I(N__22582));
    InMux I__2948 (
            .O(N__22628),
            .I(N__22582));
    InMux I__2947 (
            .O(N__22627),
            .I(N__22582));
    InMux I__2946 (
            .O(N__22626),
            .I(N__22582));
    InMux I__2945 (
            .O(N__22625),
            .I(N__22582));
    InMux I__2944 (
            .O(N__22624),
            .I(N__22582));
    InMux I__2943 (
            .O(N__22621),
            .I(N__22577));
    InMux I__2942 (
            .O(N__22618),
            .I(N__22577));
    InMux I__2941 (
            .O(N__22617),
            .I(N__22566));
    InMux I__2940 (
            .O(N__22616),
            .I(N__22566));
    InMux I__2939 (
            .O(N__22615),
            .I(N__22566));
    InMux I__2938 (
            .O(N__22614),
            .I(N__22566));
    InMux I__2937 (
            .O(N__22613),
            .I(N__22566));
    InMux I__2936 (
            .O(N__22612),
            .I(N__22561));
    InMux I__2935 (
            .O(N__22611),
            .I(N__22556));
    InMux I__2934 (
            .O(N__22610),
            .I(N__22556));
    InMux I__2933 (
            .O(N__22609),
            .I(N__22553));
    CascadeMux I__2932 (
            .O(N__22608),
            .I(N__22548));
    CascadeMux I__2931 (
            .O(N__22607),
            .I(N__22545));
    CascadeMux I__2930 (
            .O(N__22606),
            .I(N__22542));
    InMux I__2929 (
            .O(N__22603),
            .I(N__22538));
    InMux I__2928 (
            .O(N__22602),
            .I(N__22533));
    InMux I__2927 (
            .O(N__22599),
            .I(N__22533));
    InMux I__2926 (
            .O(N__22598),
            .I(N__22528));
    InMux I__2925 (
            .O(N__22597),
            .I(N__22528));
    LocalMux I__2924 (
            .O(N__22582),
            .I(N__22525));
    LocalMux I__2923 (
            .O(N__22577),
            .I(N__22520));
    LocalMux I__2922 (
            .O(N__22566),
            .I(N__22520));
    InMux I__2921 (
            .O(N__22565),
            .I(N__22515));
    InMux I__2920 (
            .O(N__22564),
            .I(N__22515));
    LocalMux I__2919 (
            .O(N__22561),
            .I(N__22510));
    LocalMux I__2918 (
            .O(N__22556),
            .I(N__22510));
    LocalMux I__2917 (
            .O(N__22553),
            .I(N__22507));
    InMux I__2916 (
            .O(N__22552),
            .I(N__22494));
    InMux I__2915 (
            .O(N__22551),
            .I(N__22494));
    InMux I__2914 (
            .O(N__22548),
            .I(N__22494));
    InMux I__2913 (
            .O(N__22545),
            .I(N__22494));
    InMux I__2912 (
            .O(N__22542),
            .I(N__22494));
    InMux I__2911 (
            .O(N__22541),
            .I(N__22494));
    LocalMux I__2910 (
            .O(N__22538),
            .I(N__22491));
    LocalMux I__2909 (
            .O(N__22533),
            .I(N__22488));
    LocalMux I__2908 (
            .O(N__22528),
            .I(N__22485));
    Span4Mux_h I__2907 (
            .O(N__22525),
            .I(N__22482));
    Span4Mux_h I__2906 (
            .O(N__22520),
            .I(N__22479));
    LocalMux I__2905 (
            .O(N__22515),
            .I(N__22472));
    Span4Mux_v I__2904 (
            .O(N__22510),
            .I(N__22472));
    Span4Mux_h I__2903 (
            .O(N__22507),
            .I(N__22472));
    LocalMux I__2902 (
            .O(N__22494),
            .I(N__22465));
    Span12Mux_v I__2901 (
            .O(N__22491),
            .I(N__22465));
    Span12Mux_v I__2900 (
            .O(N__22488),
            .I(N__22465));
    Odrv12 I__2899 (
            .O(N__22485),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2898 (
            .O(N__22482),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2897 (
            .O(N__22479),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv4 I__2896 (
            .O(N__22472),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    Odrv12 I__2895 (
            .O(N__22465),
            .I(\current_shift_inst.PI_CTRL.N_46 ));
    InMux I__2894 (
            .O(N__22454),
            .I(N__22451));
    LocalMux I__2893 (
            .O(N__22451),
            .I(N__22448));
    Odrv12 I__2892 (
            .O(N__22448),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__2891 (
            .O(N__22445),
            .I(N__22442));
    LocalMux I__2890 (
            .O(N__22442),
            .I(N__22439));
    Odrv4 I__2889 (
            .O(N__22439),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__2888 (
            .O(N__22436),
            .I(N__22430));
    InMux I__2887 (
            .O(N__22435),
            .I(N__22430));
    LocalMux I__2886 (
            .O(N__22430),
            .I(N__22427));
    Odrv4 I__2885 (
            .O(N__22427),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    CascadeMux I__2884 (
            .O(N__22424),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16_cascade_ ));
    InMux I__2883 (
            .O(N__22421),
            .I(N__22417));
    InMux I__2882 (
            .O(N__22420),
            .I(N__22414));
    LocalMux I__2881 (
            .O(N__22417),
            .I(N__22411));
    LocalMux I__2880 (
            .O(N__22414),
            .I(N__22408));
    Span4Mux_v I__2879 (
            .O(N__22411),
            .I(N__22405));
    Odrv4 I__2878 (
            .O(N__22408),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    Odrv4 I__2877 (
            .O(N__22405),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    InMux I__2876 (
            .O(N__22400),
            .I(N__22396));
    InMux I__2875 (
            .O(N__22399),
            .I(N__22393));
    LocalMux I__2874 (
            .O(N__22396),
            .I(N__22390));
    LocalMux I__2873 (
            .O(N__22393),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    Odrv4 I__2872 (
            .O(N__22390),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    CascadeMux I__2871 (
            .O(N__22385),
            .I(N__22381));
    InMux I__2870 (
            .O(N__22384),
            .I(N__22378));
    InMux I__2869 (
            .O(N__22381),
            .I(N__22375));
    LocalMux I__2868 (
            .O(N__22378),
            .I(N__22372));
    LocalMux I__2867 (
            .O(N__22375),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    Odrv4 I__2866 (
            .O(N__22372),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    CascadeMux I__2865 (
            .O(N__22367),
            .I(N__22364));
    InMux I__2864 (
            .O(N__22364),
            .I(N__22360));
    InMux I__2863 (
            .O(N__22363),
            .I(N__22357));
    LocalMux I__2862 (
            .O(N__22360),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__2861 (
            .O(N__22357),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    CascadeMux I__2860 (
            .O(N__22352),
            .I(N__22349));
    InMux I__2859 (
            .O(N__22349),
            .I(N__22346));
    LocalMux I__2858 (
            .O(N__22346),
            .I(N__22343));
    Span12Mux_h I__2857 (
            .O(N__22343),
            .I(N__22340));
    Odrv12 I__2856 (
            .O(N__22340),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__2855 (
            .O(N__22337),
            .I(N__22334));
    LocalMux I__2854 (
            .O(N__22334),
            .I(N__22331));
    Odrv4 I__2853 (
            .O(N__22331),
            .I(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ));
    InMux I__2852 (
            .O(N__22328),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    CascadeMux I__2851 (
            .O(N__22325),
            .I(N__22322));
    InMux I__2850 (
            .O(N__22322),
            .I(N__22319));
    LocalMux I__2849 (
            .O(N__22319),
            .I(N__22316));
    Odrv4 I__2848 (
            .O(N__22316),
            .I(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ));
    InMux I__2847 (
            .O(N__22313),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__2846 (
            .O(N__22310),
            .I(N__22307));
    LocalMux I__2845 (
            .O(N__22307),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__2844 (
            .O(N__22304),
            .I(bfn_4_25_0_));
    CascadeMux I__2843 (
            .O(N__22301),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_ ));
    CascadeMux I__2842 (
            .O(N__22298),
            .I(N__22295));
    InMux I__2841 (
            .O(N__22295),
            .I(N__22292));
    LocalMux I__2840 (
            .O(N__22292),
            .I(N__22288));
    InMux I__2839 (
            .O(N__22291),
            .I(N__22285));
    Span4Mux_v I__2838 (
            .O(N__22288),
            .I(N__22280));
    LocalMux I__2837 (
            .O(N__22285),
            .I(N__22280));
    Span4Mux_h I__2836 (
            .O(N__22280),
            .I(N__22277));
    Odrv4 I__2835 (
            .O(N__22277),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__2834 (
            .O(N__22274),
            .I(N__22271));
    LocalMux I__2833 (
            .O(N__22271),
            .I(N__22268));
    Span4Mux_h I__2832 (
            .O(N__22268),
            .I(N__22265));
    Odrv4 I__2831 (
            .O(N__22265),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    CascadeMux I__2830 (
            .O(N__22262),
            .I(N__22259));
    InMux I__2829 (
            .O(N__22259),
            .I(N__22256));
    LocalMux I__2828 (
            .O(N__22256),
            .I(N__22253));
    Span12Mux_h I__2827 (
            .O(N__22253),
            .I(N__22250));
    Odrv12 I__2826 (
            .O(N__22250),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    CascadeMux I__2825 (
            .O(N__22247),
            .I(N__22244));
    InMux I__2824 (
            .O(N__22244),
            .I(N__22241));
    LocalMux I__2823 (
            .O(N__22241),
            .I(N__22238));
    Odrv4 I__2822 (
            .O(N__22238),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ));
    InMux I__2821 (
            .O(N__22235),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__2820 (
            .O(N__22232),
            .I(N__22229));
    LocalMux I__2819 (
            .O(N__22229),
            .I(N__22226));
    Span12Mux_s9_h I__2818 (
            .O(N__22226),
            .I(N__22223));
    Span12Mux_h I__2817 (
            .O(N__22223),
            .I(N__22220));
    Odrv12 I__2816 (
            .O(N__22220),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    CascadeMux I__2815 (
            .O(N__22217),
            .I(N__22214));
    InMux I__2814 (
            .O(N__22214),
            .I(N__22211));
    LocalMux I__2813 (
            .O(N__22211),
            .I(N__22208));
    Span4Mux_h I__2812 (
            .O(N__22208),
            .I(N__22205));
    Odrv4 I__2811 (
            .O(N__22205),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    InMux I__2810 (
            .O(N__22202),
            .I(N__22199));
    LocalMux I__2809 (
            .O(N__22199),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ));
    InMux I__2808 (
            .O(N__22196),
            .I(bfn_4_24_0_));
    InMux I__2807 (
            .O(N__22193),
            .I(N__22190));
    LocalMux I__2806 (
            .O(N__22190),
            .I(N__22187));
    Span4Mux_h I__2805 (
            .O(N__22187),
            .I(N__22184));
    Sp12to4 I__2804 (
            .O(N__22184),
            .I(N__22181));
    Span12Mux_h I__2803 (
            .O(N__22181),
            .I(N__22178));
    Odrv12 I__2802 (
            .O(N__22178),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    CascadeMux I__2801 (
            .O(N__22175),
            .I(N__22172));
    InMux I__2800 (
            .O(N__22172),
            .I(N__22169));
    LocalMux I__2799 (
            .O(N__22169),
            .I(N__22166));
    Span4Mux_v I__2798 (
            .O(N__22166),
            .I(N__22163));
    Odrv4 I__2797 (
            .O(N__22163),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    InMux I__2796 (
            .O(N__22160),
            .I(N__22157));
    LocalMux I__2795 (
            .O(N__22157),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ));
    InMux I__2794 (
            .O(N__22154),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    InMux I__2793 (
            .O(N__22151),
            .I(N__22148));
    LocalMux I__2792 (
            .O(N__22148),
            .I(N__22145));
    Span12Mux_s7_h I__2791 (
            .O(N__22145),
            .I(N__22142));
    Span12Mux_h I__2790 (
            .O(N__22142),
            .I(N__22139));
    Odrv12 I__2789 (
            .O(N__22139),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__2788 (
            .O(N__22136),
            .I(N__22133));
    LocalMux I__2787 (
            .O(N__22133),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ));
    InMux I__2786 (
            .O(N__22130),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    InMux I__2785 (
            .O(N__22127),
            .I(N__22124));
    LocalMux I__2784 (
            .O(N__22124),
            .I(N__22121));
    Span12Mux_s6_h I__2783 (
            .O(N__22121),
            .I(N__22118));
    Span12Mux_h I__2782 (
            .O(N__22118),
            .I(N__22115));
    Odrv12 I__2781 (
            .O(N__22115),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__2780 (
            .O(N__22112),
            .I(N__22109));
    LocalMux I__2779 (
            .O(N__22109),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ));
    InMux I__2778 (
            .O(N__22106),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    InMux I__2777 (
            .O(N__22103),
            .I(N__22100));
    LocalMux I__2776 (
            .O(N__22100),
            .I(N__22097));
    Sp12to4 I__2775 (
            .O(N__22097),
            .I(N__22094));
    Span12Mux_h I__2774 (
            .O(N__22094),
            .I(N__22091));
    Odrv12 I__2773 (
            .O(N__22091),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__2772 (
            .O(N__22088),
            .I(N__22085));
    LocalMux I__2771 (
            .O(N__22085),
            .I(N__22082));
    Odrv4 I__2770 (
            .O(N__22082),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ));
    InMux I__2769 (
            .O(N__22079),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    InMux I__2768 (
            .O(N__22076),
            .I(N__22073));
    LocalMux I__2767 (
            .O(N__22073),
            .I(N__22070));
    Span12Mux_h I__2766 (
            .O(N__22070),
            .I(N__22067));
    Odrv12 I__2765 (
            .O(N__22067),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    CascadeMux I__2764 (
            .O(N__22064),
            .I(N__22061));
    InMux I__2763 (
            .O(N__22061),
            .I(N__22058));
    LocalMux I__2762 (
            .O(N__22058),
            .I(N__22055));
    Odrv4 I__2761 (
            .O(N__22055),
            .I(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ));
    InMux I__2760 (
            .O(N__22052),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    CascadeMux I__2759 (
            .O(N__22049),
            .I(N__22038));
    CascadeMux I__2758 (
            .O(N__22048),
            .I(N__22034));
    CascadeMux I__2757 (
            .O(N__22047),
            .I(N__22030));
    CascadeMux I__2756 (
            .O(N__22046),
            .I(N__22026));
    CascadeMux I__2755 (
            .O(N__22045),
            .I(N__22022));
    CascadeMux I__2754 (
            .O(N__22044),
            .I(N__22018));
    CascadeMux I__2753 (
            .O(N__22043),
            .I(N__22014));
    CascadeMux I__2752 (
            .O(N__22042),
            .I(N__22009));
    InMux I__2751 (
            .O(N__22041),
            .I(N__21993));
    InMux I__2750 (
            .O(N__22038),
            .I(N__21993));
    InMux I__2749 (
            .O(N__22037),
            .I(N__21993));
    InMux I__2748 (
            .O(N__22034),
            .I(N__21993));
    InMux I__2747 (
            .O(N__22033),
            .I(N__21993));
    InMux I__2746 (
            .O(N__22030),
            .I(N__21993));
    InMux I__2745 (
            .O(N__22029),
            .I(N__21993));
    InMux I__2744 (
            .O(N__22026),
            .I(N__21976));
    InMux I__2743 (
            .O(N__22025),
            .I(N__21976));
    InMux I__2742 (
            .O(N__22022),
            .I(N__21976));
    InMux I__2741 (
            .O(N__22021),
            .I(N__21976));
    InMux I__2740 (
            .O(N__22018),
            .I(N__21976));
    InMux I__2739 (
            .O(N__22017),
            .I(N__21976));
    InMux I__2738 (
            .O(N__22014),
            .I(N__21976));
    InMux I__2737 (
            .O(N__22013),
            .I(N__21976));
    InMux I__2736 (
            .O(N__22012),
            .I(N__21969));
    InMux I__2735 (
            .O(N__22009),
            .I(N__21969));
    InMux I__2734 (
            .O(N__22008),
            .I(N__21969));
    LocalMux I__2733 (
            .O(N__21993),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    LocalMux I__2732 (
            .O(N__21976),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    LocalMux I__2731 (
            .O(N__21969),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__2730 (
            .O(N__21962),
            .I(N__21959));
    LocalMux I__2729 (
            .O(N__21959),
            .I(N__21956));
    Span12Mux_s9_h I__2728 (
            .O(N__21956),
            .I(N__21953));
    Span12Mux_h I__2727 (
            .O(N__21953),
            .I(N__21950));
    Odrv12 I__2726 (
            .O(N__21950),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__2725 (
            .O(N__21947),
            .I(N__21944));
    InMux I__2724 (
            .O(N__21944),
            .I(N__21941));
    LocalMux I__2723 (
            .O(N__21941),
            .I(N__21938));
    Span4Mux_h I__2722 (
            .O(N__21938),
            .I(N__21935));
    Odrv4 I__2721 (
            .O(N__21935),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__2720 (
            .O(N__21932),
            .I(N__21929));
    LocalMux I__2719 (
            .O(N__21929),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__2718 (
            .O(N__21926),
            .I(N__21923));
    LocalMux I__2717 (
            .O(N__21923),
            .I(N__21920));
    Span4Mux_h I__2716 (
            .O(N__21920),
            .I(N__21917));
    Sp12to4 I__2715 (
            .O(N__21917),
            .I(N__21914));
    Span12Mux_h I__2714 (
            .O(N__21914),
            .I(N__21911));
    Odrv12 I__2713 (
            .O(N__21911),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__2712 (
            .O(N__21908),
            .I(N__21905));
    InMux I__2711 (
            .O(N__21905),
            .I(N__21902));
    LocalMux I__2710 (
            .O(N__21902),
            .I(N__21899));
    Span4Mux_h I__2709 (
            .O(N__21899),
            .I(N__21896));
    Odrv4 I__2708 (
            .O(N__21896),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    CascadeMux I__2707 (
            .O(N__21893),
            .I(N__21890));
    InMux I__2706 (
            .O(N__21890),
            .I(N__21887));
    LocalMux I__2705 (
            .O(N__21887),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ));
    InMux I__2704 (
            .O(N__21884),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__2703 (
            .O(N__21881),
            .I(N__21878));
    LocalMux I__2702 (
            .O(N__21878),
            .I(N__21875));
    Span12Mux_s7_h I__2701 (
            .O(N__21875),
            .I(N__21872));
    Span12Mux_h I__2700 (
            .O(N__21872),
            .I(N__21869));
    Odrv12 I__2699 (
            .O(N__21869),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__2698 (
            .O(N__21866),
            .I(N__21863));
    InMux I__2697 (
            .O(N__21863),
            .I(N__21860));
    LocalMux I__2696 (
            .O(N__21860),
            .I(N__21857));
    Span4Mux_h I__2695 (
            .O(N__21857),
            .I(N__21854));
    Odrv4 I__2694 (
            .O(N__21854),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__2693 (
            .O(N__21851),
            .I(N__21848));
    LocalMux I__2692 (
            .O(N__21848),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ));
    InMux I__2691 (
            .O(N__21845),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__2690 (
            .O(N__21842),
            .I(N__21839));
    LocalMux I__2689 (
            .O(N__21839),
            .I(N__21836));
    Span12Mux_s6_h I__2688 (
            .O(N__21836),
            .I(N__21833));
    Span12Mux_h I__2687 (
            .O(N__21833),
            .I(N__21830));
    Odrv12 I__2686 (
            .O(N__21830),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__2685 (
            .O(N__21827),
            .I(N__21824));
    InMux I__2684 (
            .O(N__21824),
            .I(N__21821));
    LocalMux I__2683 (
            .O(N__21821),
            .I(N__21818));
    Span4Mux_v I__2682 (
            .O(N__21818),
            .I(N__21815));
    Odrv4 I__2681 (
            .O(N__21815),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    CascadeMux I__2680 (
            .O(N__21812),
            .I(N__21809));
    InMux I__2679 (
            .O(N__21809),
            .I(N__21806));
    LocalMux I__2678 (
            .O(N__21806),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ));
    InMux I__2677 (
            .O(N__21803),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__2676 (
            .O(N__21800),
            .I(N__21797));
    LocalMux I__2675 (
            .O(N__21797),
            .I(N__21794));
    Span4Mux_v I__2674 (
            .O(N__21794),
            .I(N__21791));
    Odrv4 I__2673 (
            .O(N__21791),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    CascadeMux I__2672 (
            .O(N__21788),
            .I(N__21785));
    InMux I__2671 (
            .O(N__21785),
            .I(N__21782));
    LocalMux I__2670 (
            .O(N__21782),
            .I(N__21779));
    Span12Mux_s5_h I__2669 (
            .O(N__21779),
            .I(N__21776));
    Span12Mux_h I__2668 (
            .O(N__21776),
            .I(N__21773));
    Odrv12 I__2667 (
            .O(N__21773),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    InMux I__2666 (
            .O(N__21770),
            .I(N__21767));
    LocalMux I__2665 (
            .O(N__21767),
            .I(N__21764));
    Odrv4 I__2664 (
            .O(N__21764),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ));
    InMux I__2663 (
            .O(N__21761),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__2662 (
            .O(N__21758),
            .I(N__21755));
    LocalMux I__2661 (
            .O(N__21755),
            .I(N__21752));
    Span4Mux_h I__2660 (
            .O(N__21752),
            .I(N__21749));
    Odrv4 I__2659 (
            .O(N__21749),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    CascadeMux I__2658 (
            .O(N__21746),
            .I(N__21743));
    InMux I__2657 (
            .O(N__21743),
            .I(N__21740));
    LocalMux I__2656 (
            .O(N__21740),
            .I(N__21737));
    Span12Mux_h I__2655 (
            .O(N__21737),
            .I(N__21734));
    Odrv12 I__2654 (
            .O(N__21734),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__2653 (
            .O(N__21731),
            .I(N__21728));
    InMux I__2652 (
            .O(N__21728),
            .I(N__21725));
    LocalMux I__2651 (
            .O(N__21725),
            .I(N__21722));
    Odrv4 I__2650 (
            .O(N__21722),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ));
    InMux I__2649 (
            .O(N__21719),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__2648 (
            .O(N__21716),
            .I(N__21713));
    LocalMux I__2647 (
            .O(N__21713),
            .I(N__21710));
    Span4Mux_h I__2646 (
            .O(N__21710),
            .I(N__21707));
    Odrv4 I__2645 (
            .O(N__21707),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    CascadeMux I__2644 (
            .O(N__21704),
            .I(N__21701));
    InMux I__2643 (
            .O(N__21701),
            .I(N__21698));
    LocalMux I__2642 (
            .O(N__21698),
            .I(N__21695));
    Span12Mux_h I__2641 (
            .O(N__21695),
            .I(N__21692));
    Odrv12 I__2640 (
            .O(N__21692),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    InMux I__2639 (
            .O(N__21689),
            .I(N__21686));
    LocalMux I__2638 (
            .O(N__21686),
            .I(N__21683));
    Odrv4 I__2637 (
            .O(N__21683),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ));
    InMux I__2636 (
            .O(N__21680),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    CascadeMux I__2635 (
            .O(N__21677),
            .I(N__21674));
    InMux I__2634 (
            .O(N__21674),
            .I(N__21671));
    LocalMux I__2633 (
            .O(N__21671),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    InMux I__2632 (
            .O(N__21668),
            .I(N__21665));
    LocalMux I__2631 (
            .O(N__21665),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__2630 (
            .O(N__21662),
            .I(N__21659));
    LocalMux I__2629 (
            .O(N__21659),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    InMux I__2628 (
            .O(N__21656),
            .I(N__21653));
    LocalMux I__2627 (
            .O(N__21653),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__2626 (
            .O(N__21650),
            .I(N__21647));
    LocalMux I__2625 (
            .O(N__21647),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__2624 (
            .O(N__21644),
            .I(N__21641));
    LocalMux I__2623 (
            .O(N__21641),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__2622 (
            .O(N__21638),
            .I(N__21634));
    InMux I__2621 (
            .O(N__21637),
            .I(N__21631));
    LocalMux I__2620 (
            .O(N__21634),
            .I(N__21628));
    LocalMux I__2619 (
            .O(N__21631),
            .I(N__21625));
    Span4Mux_h I__2618 (
            .O(N__21628),
            .I(N__21622));
    Odrv4 I__2617 (
            .O(N__21625),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    Odrv4 I__2616 (
            .O(N__21622),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__2615 (
            .O(N__21617),
            .I(N__21614));
    LocalMux I__2614 (
            .O(N__21614),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    InMux I__2613 (
            .O(N__21611),
            .I(N__21608));
    LocalMux I__2612 (
            .O(N__21608),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__2611 (
            .O(N__21605),
            .I(N__21602));
    LocalMux I__2610 (
            .O(N__21602),
            .I(N__21599));
    Span4Mux_v I__2609 (
            .O(N__21599),
            .I(N__21593));
    InMux I__2608 (
            .O(N__21598),
            .I(N__21590));
    InMux I__2607 (
            .O(N__21597),
            .I(N__21587));
    InMux I__2606 (
            .O(N__21596),
            .I(N__21584));
    Odrv4 I__2605 (
            .O(N__21593),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__2604 (
            .O(N__21590),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__2603 (
            .O(N__21587),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__2602 (
            .O(N__21584),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__2601 (
            .O(N__21575),
            .I(N__21571));
    CascadeMux I__2600 (
            .O(N__21574),
            .I(N__21567));
    LocalMux I__2599 (
            .O(N__21571),
            .I(N__21563));
    InMux I__2598 (
            .O(N__21570),
            .I(N__21560));
    InMux I__2597 (
            .O(N__21567),
            .I(N__21557));
    InMux I__2596 (
            .O(N__21566),
            .I(N__21554));
    Odrv12 I__2595 (
            .O(N__21563),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__2594 (
            .O(N__21560),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__2593 (
            .O(N__21557),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__2592 (
            .O(N__21554),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__2591 (
            .O(N__21545),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ));
    InMux I__2590 (
            .O(N__21542),
            .I(N__21539));
    LocalMux I__2589 (
            .O(N__21539),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    CascadeMux I__2588 (
            .O(N__21536),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ));
    InMux I__2587 (
            .O(N__21533),
            .I(N__21530));
    LocalMux I__2586 (
            .O(N__21530),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    InMux I__2585 (
            .O(N__21527),
            .I(N__21524));
    LocalMux I__2584 (
            .O(N__21524),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__2583 (
            .O(N__21521),
            .I(N__21518));
    LocalMux I__2582 (
            .O(N__21518),
            .I(N__21512));
    InMux I__2581 (
            .O(N__21517),
            .I(N__21509));
    InMux I__2580 (
            .O(N__21516),
            .I(N__21504));
    InMux I__2579 (
            .O(N__21515),
            .I(N__21504));
    Odrv12 I__2578 (
            .O(N__21512),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__2577 (
            .O(N__21509),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__2576 (
            .O(N__21504),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__2575 (
            .O(N__21497),
            .I(N__21494));
    LocalMux I__2574 (
            .O(N__21494),
            .I(N__21488));
    InMux I__2573 (
            .O(N__21493),
            .I(N__21485));
    InMux I__2572 (
            .O(N__21492),
            .I(N__21480));
    InMux I__2571 (
            .O(N__21491),
            .I(N__21480));
    Odrv12 I__2570 (
            .O(N__21488),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__2569 (
            .O(N__21485),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__2568 (
            .O(N__21480),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    CascadeMux I__2567 (
            .O(N__21473),
            .I(N__21470));
    InMux I__2566 (
            .O(N__21470),
            .I(N__21467));
    LocalMux I__2565 (
            .O(N__21467),
            .I(N__21463));
    CascadeMux I__2564 (
            .O(N__21466),
            .I(N__21459));
    Span4Mux_v I__2563 (
            .O(N__21463),
            .I(N__21455));
    InMux I__2562 (
            .O(N__21462),
            .I(N__21452));
    InMux I__2561 (
            .O(N__21459),
            .I(N__21447));
    InMux I__2560 (
            .O(N__21458),
            .I(N__21447));
    Odrv4 I__2559 (
            .O(N__21455),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__2558 (
            .O(N__21452),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__2557 (
            .O(N__21447),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    CascadeMux I__2556 (
            .O(N__21440),
            .I(N__21436));
    CascadeMux I__2555 (
            .O(N__21439),
            .I(N__21432));
    InMux I__2554 (
            .O(N__21436),
            .I(N__21429));
    InMux I__2553 (
            .O(N__21435),
            .I(N__21424));
    InMux I__2552 (
            .O(N__21432),
            .I(N__21424));
    LocalMux I__2551 (
            .O(N__21429),
            .I(N__21420));
    LocalMux I__2550 (
            .O(N__21424),
            .I(N__21417));
    InMux I__2549 (
            .O(N__21423),
            .I(N__21414));
    Span4Mux_v I__2548 (
            .O(N__21420),
            .I(N__21409));
    Span4Mux_h I__2547 (
            .O(N__21417),
            .I(N__21409));
    LocalMux I__2546 (
            .O(N__21414),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__2545 (
            .O(N__21409),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    CascadeMux I__2544 (
            .O(N__21404),
            .I(N__21401));
    InMux I__2543 (
            .O(N__21401),
            .I(N__21398));
    LocalMux I__2542 (
            .O(N__21398),
            .I(N__21393));
    InMux I__2541 (
            .O(N__21397),
            .I(N__21390));
    InMux I__2540 (
            .O(N__21396),
            .I(N__21386));
    Span4Mux_v I__2539 (
            .O(N__21393),
            .I(N__21381));
    LocalMux I__2538 (
            .O(N__21390),
            .I(N__21381));
    InMux I__2537 (
            .O(N__21389),
            .I(N__21378));
    LocalMux I__2536 (
            .O(N__21386),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    Odrv4 I__2535 (
            .O(N__21381),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__2534 (
            .O(N__21378),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    CascadeMux I__2533 (
            .O(N__21371),
            .I(N__21368));
    InMux I__2532 (
            .O(N__21368),
            .I(N__21365));
    LocalMux I__2531 (
            .O(N__21365),
            .I(N__21360));
    InMux I__2530 (
            .O(N__21364),
            .I(N__21357));
    InMux I__2529 (
            .O(N__21363),
            .I(N__21353));
    Span4Mux_v I__2528 (
            .O(N__21360),
            .I(N__21348));
    LocalMux I__2527 (
            .O(N__21357),
            .I(N__21348));
    InMux I__2526 (
            .O(N__21356),
            .I(N__21345));
    LocalMux I__2525 (
            .O(N__21353),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__2524 (
            .O(N__21348),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__2523 (
            .O(N__21345),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__2522 (
            .O(N__21338),
            .I(N__21335));
    LocalMux I__2521 (
            .O(N__21335),
            .I(N__21329));
    InMux I__2520 (
            .O(N__21334),
            .I(N__21326));
    InMux I__2519 (
            .O(N__21333),
            .I(N__21321));
    InMux I__2518 (
            .O(N__21332),
            .I(N__21321));
    Odrv12 I__2517 (
            .O(N__21329),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__2516 (
            .O(N__21326),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__2515 (
            .O(N__21321),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__2514 (
            .O(N__21314),
            .I(N__21310));
    CascadeMux I__2513 (
            .O(N__21313),
            .I(N__21306));
    InMux I__2512 (
            .O(N__21310),
            .I(N__21303));
    InMux I__2511 (
            .O(N__21309),
            .I(N__21300));
    InMux I__2510 (
            .O(N__21306),
            .I(N__21297));
    LocalMux I__2509 (
            .O(N__21303),
            .I(N__21293));
    LocalMux I__2508 (
            .O(N__21300),
            .I(N__21288));
    LocalMux I__2507 (
            .O(N__21297),
            .I(N__21288));
    InMux I__2506 (
            .O(N__21296),
            .I(N__21285));
    Span4Mux_v I__2505 (
            .O(N__21293),
            .I(N__21280));
    Span4Mux_v I__2504 (
            .O(N__21288),
            .I(N__21280));
    LocalMux I__2503 (
            .O(N__21285),
            .I(N__21277));
    Odrv4 I__2502 (
            .O(N__21280),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__2501 (
            .O(N__21277),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__2500 (
            .O(N__21272),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ));
    InMux I__2499 (
            .O(N__21269),
            .I(N__21266));
    LocalMux I__2498 (
            .O(N__21266),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ));
    InMux I__2497 (
            .O(N__21263),
            .I(N__21260));
    LocalMux I__2496 (
            .O(N__21260),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__2495 (
            .O(N__21257),
            .I(N__21254));
    LocalMux I__2494 (
            .O(N__21254),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    CascadeMux I__2493 (
            .O(N__21251),
            .I(N__21248));
    InMux I__2492 (
            .O(N__21248),
            .I(N__21245));
    LocalMux I__2491 (
            .O(N__21245),
            .I(N__21241));
    InMux I__2490 (
            .O(N__21244),
            .I(N__21236));
    Span4Mux_v I__2489 (
            .O(N__21241),
            .I(N__21233));
    InMux I__2488 (
            .O(N__21240),
            .I(N__21228));
    InMux I__2487 (
            .O(N__21239),
            .I(N__21228));
    LocalMux I__2486 (
            .O(N__21236),
            .I(N__21225));
    Odrv4 I__2485 (
            .O(N__21233),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__2484 (
            .O(N__21228),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__2483 (
            .O(N__21225),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    InMux I__2482 (
            .O(N__21218),
            .I(N__21215));
    LocalMux I__2481 (
            .O(N__21215),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ));
    InMux I__2480 (
            .O(N__21212),
            .I(N__21209));
    LocalMux I__2479 (
            .O(N__21209),
            .I(N__21206));
    Odrv12 I__2478 (
            .O(N__21206),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    InMux I__2477 (
            .O(N__21203),
            .I(N__21200));
    LocalMux I__2476 (
            .O(N__21200),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    CascadeMux I__2475 (
            .O(N__21197),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ));
    InMux I__2474 (
            .O(N__21194),
            .I(N__21191));
    LocalMux I__2473 (
            .O(N__21191),
            .I(N__21188));
    Span4Mux_v I__2472 (
            .O(N__21188),
            .I(N__21182));
    InMux I__2471 (
            .O(N__21187),
            .I(N__21179));
    InMux I__2470 (
            .O(N__21186),
            .I(N__21174));
    InMux I__2469 (
            .O(N__21185),
            .I(N__21174));
    Odrv4 I__2468 (
            .O(N__21182),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__2467 (
            .O(N__21179),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__2466 (
            .O(N__21174),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__2465 (
            .O(N__21167),
            .I(N__21164));
    InMux I__2464 (
            .O(N__21164),
            .I(N__21161));
    LocalMux I__2463 (
            .O(N__21161),
            .I(N__21158));
    Span4Mux_v I__2462 (
            .O(N__21158),
            .I(N__21152));
    InMux I__2461 (
            .O(N__21157),
            .I(N__21149));
    InMux I__2460 (
            .O(N__21156),
            .I(N__21144));
    InMux I__2459 (
            .O(N__21155),
            .I(N__21144));
    Odrv4 I__2458 (
            .O(N__21152),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__2457 (
            .O(N__21149),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    LocalMux I__2456 (
            .O(N__21144),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    CascadeMux I__2455 (
            .O(N__21137),
            .I(N__21134));
    InMux I__2454 (
            .O(N__21134),
            .I(N__21131));
    LocalMux I__2453 (
            .O(N__21131),
            .I(N__21126));
    CascadeMux I__2452 (
            .O(N__21130),
            .I(N__21123));
    CascadeMux I__2451 (
            .O(N__21129),
            .I(N__21120));
    Span4Mux_v I__2450 (
            .O(N__21126),
            .I(N__21116));
    InMux I__2449 (
            .O(N__21123),
            .I(N__21111));
    InMux I__2448 (
            .O(N__21120),
            .I(N__21111));
    InMux I__2447 (
            .O(N__21119),
            .I(N__21108));
    Odrv4 I__2446 (
            .O(N__21116),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__2445 (
            .O(N__21111),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__2444 (
            .O(N__21108),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__2443 (
            .O(N__21101),
            .I(N__21098));
    InMux I__2442 (
            .O(N__21098),
            .I(N__21095));
    LocalMux I__2441 (
            .O(N__21095),
            .I(N__21092));
    Span4Mux_v I__2440 (
            .O(N__21092),
            .I(N__21086));
    InMux I__2439 (
            .O(N__21091),
            .I(N__21083));
    InMux I__2438 (
            .O(N__21090),
            .I(N__21080));
    InMux I__2437 (
            .O(N__21089),
            .I(N__21077));
    Odrv4 I__2436 (
            .O(N__21086),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__2435 (
            .O(N__21083),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__2434 (
            .O(N__21080),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__2433 (
            .O(N__21077),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    CascadeMux I__2432 (
            .O(N__21068),
            .I(N__21065));
    InMux I__2431 (
            .O(N__21065),
            .I(N__21062));
    LocalMux I__2430 (
            .O(N__21062),
            .I(N__21056));
    InMux I__2429 (
            .O(N__21061),
            .I(N__21053));
    InMux I__2428 (
            .O(N__21060),
            .I(N__21048));
    InMux I__2427 (
            .O(N__21059),
            .I(N__21048));
    Odrv12 I__2426 (
            .O(N__21056),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__2425 (
            .O(N__21053),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__2424 (
            .O(N__21048),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    InMux I__2423 (
            .O(N__21041),
            .I(N__21038));
    LocalMux I__2422 (
            .O(N__21038),
            .I(N__21033));
    InMux I__2421 (
            .O(N__21037),
            .I(N__21027));
    InMux I__2420 (
            .O(N__21036),
            .I(N__21027));
    Span12Mux_h I__2419 (
            .O(N__21033),
            .I(N__21024));
    InMux I__2418 (
            .O(N__21032),
            .I(N__21021));
    LocalMux I__2417 (
            .O(N__21027),
            .I(N__21018));
    Odrv12 I__2416 (
            .O(N__21024),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__2415 (
            .O(N__21021),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__2414 (
            .O(N__21018),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__2413 (
            .O(N__21011),
            .I(N__21006));
    CascadeMux I__2412 (
            .O(N__21010),
            .I(N__21002));
    CascadeMux I__2411 (
            .O(N__21009),
            .I(N__20999));
    LocalMux I__2410 (
            .O(N__21006),
            .I(N__20996));
    InMux I__2409 (
            .O(N__21005),
            .I(N__20993));
    InMux I__2408 (
            .O(N__21002),
            .I(N__20988));
    InMux I__2407 (
            .O(N__20999),
            .I(N__20988));
    Odrv12 I__2406 (
            .O(N__20996),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__2405 (
            .O(N__20993),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__2404 (
            .O(N__20988),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    CascadeMux I__2403 (
            .O(N__20981),
            .I(N__20978));
    InMux I__2402 (
            .O(N__20978),
            .I(N__20975));
    LocalMux I__2401 (
            .O(N__20975),
            .I(N__20969));
    InMux I__2400 (
            .O(N__20974),
            .I(N__20966));
    InMux I__2399 (
            .O(N__20973),
            .I(N__20961));
    InMux I__2398 (
            .O(N__20972),
            .I(N__20961));
    Odrv12 I__2397 (
            .O(N__20969),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__2396 (
            .O(N__20966),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__2395 (
            .O(N__20961),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    CascadeMux I__2394 (
            .O(N__20954),
            .I(N__20951));
    InMux I__2393 (
            .O(N__20951),
            .I(N__20948));
    LocalMux I__2392 (
            .O(N__20948),
            .I(N__20942));
    InMux I__2391 (
            .O(N__20947),
            .I(N__20939));
    InMux I__2390 (
            .O(N__20946),
            .I(N__20936));
    InMux I__2389 (
            .O(N__20945),
            .I(N__20933));
    Odrv4 I__2388 (
            .O(N__20942),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__2387 (
            .O(N__20939),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__2386 (
            .O(N__20936),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__2385 (
            .O(N__20933),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__2384 (
            .O(N__20924),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__2383 (
            .O(N__20921),
            .I(N__20918));
    LocalMux I__2382 (
            .O(N__20918),
            .I(N__20915));
    Span12Mux_h I__2381 (
            .O(N__20915),
            .I(N__20912));
    Odrv12 I__2380 (
            .O(N__20912),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    CascadeMux I__2379 (
            .O(N__20909),
            .I(N__20906));
    InMux I__2378 (
            .O(N__20906),
            .I(N__20903));
    LocalMux I__2377 (
            .O(N__20903),
            .I(N__20900));
    Odrv4 I__2376 (
            .O(N__20900),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    CascadeMux I__2375 (
            .O(N__20897),
            .I(N__20894));
    InMux I__2374 (
            .O(N__20894),
            .I(N__20891));
    LocalMux I__2373 (
            .O(N__20891),
            .I(N__20888));
    Odrv12 I__2372 (
            .O(N__20888),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__2371 (
            .O(N__20885),
            .I(N__20881));
    InMux I__2370 (
            .O(N__20884),
            .I(N__20877));
    InMux I__2369 (
            .O(N__20881),
            .I(N__20874));
    InMux I__2368 (
            .O(N__20880),
            .I(N__20871));
    LocalMux I__2367 (
            .O(N__20877),
            .I(N__20868));
    LocalMux I__2366 (
            .O(N__20874),
            .I(N__20865));
    LocalMux I__2365 (
            .O(N__20871),
            .I(N__20862));
    Span4Mux_h I__2364 (
            .O(N__20868),
            .I(N__20859));
    Span4Mux_h I__2363 (
            .O(N__20865),
            .I(N__20856));
    Span4Mux_v I__2362 (
            .O(N__20862),
            .I(N__20853));
    Odrv4 I__2361 (
            .O(N__20859),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__2360 (
            .O(N__20856),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__2359 (
            .O(N__20853),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    CascadeMux I__2358 (
            .O(N__20846),
            .I(N__20842));
    InMux I__2357 (
            .O(N__20845),
            .I(N__20839));
    InMux I__2356 (
            .O(N__20842),
            .I(N__20835));
    LocalMux I__2355 (
            .O(N__20839),
            .I(N__20831));
    CascadeMux I__2354 (
            .O(N__20838),
            .I(N__20828));
    LocalMux I__2353 (
            .O(N__20835),
            .I(N__20825));
    InMux I__2352 (
            .O(N__20834),
            .I(N__20821));
    Span4Mux_v I__2351 (
            .O(N__20831),
            .I(N__20818));
    InMux I__2350 (
            .O(N__20828),
            .I(N__20815));
    Span4Mux_h I__2349 (
            .O(N__20825),
            .I(N__20812));
    InMux I__2348 (
            .O(N__20824),
            .I(N__20809));
    LocalMux I__2347 (
            .O(N__20821),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__2346 (
            .O(N__20818),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__2345 (
            .O(N__20815),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__2344 (
            .O(N__20812),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__2343 (
            .O(N__20809),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__2342 (
            .O(N__20798),
            .I(\current_shift_inst.PI_CTRL.N_77_cascade_ ));
    CascadeMux I__2341 (
            .O(N__20795),
            .I(N__20792));
    InMux I__2340 (
            .O(N__20792),
            .I(N__20788));
    InMux I__2339 (
            .O(N__20791),
            .I(N__20784));
    LocalMux I__2338 (
            .O(N__20788),
            .I(N__20781));
    InMux I__2337 (
            .O(N__20787),
            .I(N__20777));
    LocalMux I__2336 (
            .O(N__20784),
            .I(N__20774));
    Span4Mux_v I__2335 (
            .O(N__20781),
            .I(N__20771));
    InMux I__2334 (
            .O(N__20780),
            .I(N__20768));
    LocalMux I__2333 (
            .O(N__20777),
            .I(N__20765));
    Odrv4 I__2332 (
            .O(N__20774),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__2331 (
            .O(N__20771),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__2330 (
            .O(N__20768),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__2329 (
            .O(N__20765),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__2328 (
            .O(N__20756),
            .I(N__20753));
    LocalMux I__2327 (
            .O(N__20753),
            .I(N__20750));
    Odrv4 I__2326 (
            .O(N__20750),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__2325 (
            .O(N__20747),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__2324 (
            .O(N__20744),
            .I(N__20741));
    LocalMux I__2323 (
            .O(N__20741),
            .I(N__20738));
    Odrv4 I__2322 (
            .O(N__20738),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__2321 (
            .O(N__20735),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__2320 (
            .O(N__20732),
            .I(N__20729));
    LocalMux I__2319 (
            .O(N__20729),
            .I(N__20726));
    Odrv12 I__2318 (
            .O(N__20726),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__2317 (
            .O(N__20723),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__2316 (
            .O(N__20720),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    InMux I__2315 (
            .O(N__20717),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__2314 (
            .O(N__20714),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__2313 (
            .O(N__20711),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__2312 (
            .O(N__20708),
            .I(bfn_3_25_0_));
    CascadeMux I__2311 (
            .O(N__20705),
            .I(N__20701));
    InMux I__2310 (
            .O(N__20704),
            .I(N__20696));
    InMux I__2309 (
            .O(N__20701),
            .I(N__20696));
    LocalMux I__2308 (
            .O(N__20696),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2307 (
            .O(N__20693),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2306 (
            .O(N__20690),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2305 (
            .O(N__20687),
            .I(N__20683));
    CascadeMux I__2304 (
            .O(N__20686),
            .I(N__20680));
    LocalMux I__2303 (
            .O(N__20683),
            .I(N__20676));
    InMux I__2302 (
            .O(N__20680),
            .I(N__20673));
    InMux I__2301 (
            .O(N__20679),
            .I(N__20670));
    Span4Mux_v I__2300 (
            .O(N__20676),
            .I(N__20664));
    LocalMux I__2299 (
            .O(N__20673),
            .I(N__20664));
    LocalMux I__2298 (
            .O(N__20670),
            .I(N__20661));
    InMux I__2297 (
            .O(N__20669),
            .I(N__20658));
    Span4Mux_v I__2296 (
            .O(N__20664),
            .I(N__20655));
    Sp12to4 I__2295 (
            .O(N__20661),
            .I(N__20650));
    LocalMux I__2294 (
            .O(N__20658),
            .I(N__20650));
    Odrv4 I__2293 (
            .O(N__20655),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv12 I__2292 (
            .O(N__20650),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2291 (
            .O(N__20645),
            .I(N__20642));
    LocalMux I__2290 (
            .O(N__20642),
            .I(N__20638));
    InMux I__2289 (
            .O(N__20641),
            .I(N__20635));
    Span4Mux_s3_h I__2288 (
            .O(N__20638),
            .I(N__20631));
    LocalMux I__2287 (
            .O(N__20635),
            .I(N__20628));
    InMux I__2286 (
            .O(N__20634),
            .I(N__20625));
    Span4Mux_v I__2285 (
            .O(N__20631),
            .I(N__20622));
    Sp12to4 I__2284 (
            .O(N__20628),
            .I(N__20617));
    LocalMux I__2283 (
            .O(N__20625),
            .I(N__20617));
    Odrv4 I__2282 (
            .O(N__20622),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv12 I__2281 (
            .O(N__20617),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2280 (
            .O(N__20612),
            .I(N__20609));
    LocalMux I__2279 (
            .O(N__20609),
            .I(\current_shift_inst.PI_CTRL.N_98 ));
    CascadeMux I__2278 (
            .O(N__20606),
            .I(N__20603));
    InMux I__2277 (
            .O(N__20603),
            .I(N__20600));
    LocalMux I__2276 (
            .O(N__20600),
            .I(N__20596));
    InMux I__2275 (
            .O(N__20599),
            .I(N__20593));
    Span4Mux_v I__2274 (
            .O(N__20596),
            .I(N__20590));
    LocalMux I__2273 (
            .O(N__20593),
            .I(N__20587));
    Odrv4 I__2272 (
            .O(N__20590),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    Odrv4 I__2271 (
            .O(N__20587),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2270 (
            .O(N__20582),
            .I(N__20578));
    InMux I__2269 (
            .O(N__20581),
            .I(N__20575));
    LocalMux I__2268 (
            .O(N__20578),
            .I(N__20572));
    LocalMux I__2267 (
            .O(N__20575),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    Odrv4 I__2266 (
            .O(N__20572),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    CascadeMux I__2265 (
            .O(N__20567),
            .I(N__20564));
    InMux I__2264 (
            .O(N__20564),
            .I(N__20560));
    InMux I__2263 (
            .O(N__20563),
            .I(N__20557));
    LocalMux I__2262 (
            .O(N__20560),
            .I(N__20552));
    LocalMux I__2261 (
            .O(N__20557),
            .I(N__20552));
    Odrv4 I__2260 (
            .O(N__20552),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    CascadeMux I__2259 (
            .O(N__20549),
            .I(N__20545));
    InMux I__2258 (
            .O(N__20548),
            .I(N__20542));
    InMux I__2257 (
            .O(N__20545),
            .I(N__20539));
    LocalMux I__2256 (
            .O(N__20542),
            .I(N__20536));
    LocalMux I__2255 (
            .O(N__20539),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    Odrv4 I__2254 (
            .O(N__20536),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2253 (
            .O(N__20531),
            .I(N__20528));
    LocalMux I__2252 (
            .O(N__20528),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ));
    InMux I__2251 (
            .O(N__20525),
            .I(N__20521));
    InMux I__2250 (
            .O(N__20524),
            .I(N__20517));
    LocalMux I__2249 (
            .O(N__20521),
            .I(N__20514));
    InMux I__2248 (
            .O(N__20520),
            .I(N__20511));
    LocalMux I__2247 (
            .O(N__20517),
            .I(N__20508));
    Span12Mux_s3_h I__2246 (
            .O(N__20514),
            .I(N__20503));
    LocalMux I__2245 (
            .O(N__20511),
            .I(N__20503));
    Odrv4 I__2244 (
            .O(N__20508),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    Odrv12 I__2243 (
            .O(N__20503),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    CascadeMux I__2242 (
            .O(N__20498),
            .I(N__20495));
    InMux I__2241 (
            .O(N__20495),
            .I(N__20492));
    LocalMux I__2240 (
            .O(N__20492),
            .I(N__20488));
    InMux I__2239 (
            .O(N__20491),
            .I(N__20485));
    Span4Mux_s3_h I__2238 (
            .O(N__20488),
            .I(N__20481));
    LocalMux I__2237 (
            .O(N__20485),
            .I(N__20478));
    InMux I__2236 (
            .O(N__20484),
            .I(N__20475));
    Span4Mux_v I__2235 (
            .O(N__20481),
            .I(N__20472));
    Span4Mux_v I__2234 (
            .O(N__20478),
            .I(N__20467));
    LocalMux I__2233 (
            .O(N__20475),
            .I(N__20467));
    Odrv4 I__2232 (
            .O(N__20472),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv4 I__2231 (
            .O(N__20467),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2230 (
            .O(N__20462),
            .I(N__20458));
    CascadeMux I__2229 (
            .O(N__20461),
            .I(N__20454));
    LocalMux I__2228 (
            .O(N__20458),
            .I(N__20451));
    InMux I__2227 (
            .O(N__20457),
            .I(N__20448));
    InMux I__2226 (
            .O(N__20454),
            .I(N__20445));
    Span12Mux_v I__2225 (
            .O(N__20451),
            .I(N__20442));
    LocalMux I__2224 (
            .O(N__20448),
            .I(N__20439));
    LocalMux I__2223 (
            .O(N__20445),
            .I(N__20436));
    Odrv12 I__2222 (
            .O(N__20442),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv12 I__2221 (
            .O(N__20439),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv4 I__2220 (
            .O(N__20436),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2219 (
            .O(N__20429),
            .I(N__20426));
    LocalMux I__2218 (
            .O(N__20426),
            .I(N__20422));
    InMux I__2217 (
            .O(N__20425),
            .I(N__20419));
    Span4Mux_h I__2216 (
            .O(N__20422),
            .I(N__20415));
    LocalMux I__2215 (
            .O(N__20419),
            .I(N__20412));
    InMux I__2214 (
            .O(N__20418),
            .I(N__20409));
    Span4Mux_v I__2213 (
            .O(N__20415),
            .I(N__20406));
    Span4Mux_v I__2212 (
            .O(N__20412),
            .I(N__20401));
    LocalMux I__2211 (
            .O(N__20409),
            .I(N__20401));
    Odrv4 I__2210 (
            .O(N__20406),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2209 (
            .O(N__20401),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    CascadeMux I__2208 (
            .O(N__20396),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ));
    InMux I__2207 (
            .O(N__20393),
            .I(N__20390));
    LocalMux I__2206 (
            .O(N__20390),
            .I(N__20387));
    Span4Mux_s3_h I__2205 (
            .O(N__20387),
            .I(N__20383));
    InMux I__2204 (
            .O(N__20386),
            .I(N__20380));
    Span4Mux_v I__2203 (
            .O(N__20383),
            .I(N__20376));
    LocalMux I__2202 (
            .O(N__20380),
            .I(N__20373));
    InMux I__2201 (
            .O(N__20379),
            .I(N__20370));
    Odrv4 I__2200 (
            .O(N__20376),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv12 I__2199 (
            .O(N__20373),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    LocalMux I__2198 (
            .O(N__20370),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    CascadeMux I__2197 (
            .O(N__20363),
            .I(N__20360));
    InMux I__2196 (
            .O(N__20360),
            .I(N__20357));
    LocalMux I__2195 (
            .O(N__20357),
            .I(N__20353));
    CascadeMux I__2194 (
            .O(N__20356),
            .I(N__20350));
    Span4Mux_v I__2193 (
            .O(N__20353),
            .I(N__20347));
    InMux I__2192 (
            .O(N__20350),
            .I(N__20344));
    Odrv4 I__2191 (
            .O(N__20347),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__2190 (
            .O(N__20344),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    InMux I__2189 (
            .O(N__20339),
            .I(N__20335));
    InMux I__2188 (
            .O(N__20338),
            .I(N__20332));
    LocalMux I__2187 (
            .O(N__20335),
            .I(N__20329));
    LocalMux I__2186 (
            .O(N__20332),
            .I(N__20325));
    Span4Mux_h I__2185 (
            .O(N__20329),
            .I(N__20322));
    InMux I__2184 (
            .O(N__20328),
            .I(N__20319));
    Span4Mux_s1_h I__2183 (
            .O(N__20325),
            .I(N__20316));
    Odrv4 I__2182 (
            .O(N__20322),
            .I(pwm_duty_input_3));
    LocalMux I__2181 (
            .O(N__20319),
            .I(pwm_duty_input_3));
    Odrv4 I__2180 (
            .O(N__20316),
            .I(pwm_duty_input_3));
    InMux I__2179 (
            .O(N__20309),
            .I(N__20305));
    InMux I__2178 (
            .O(N__20308),
            .I(N__20301));
    LocalMux I__2177 (
            .O(N__20305),
            .I(N__20298));
    InMux I__2176 (
            .O(N__20304),
            .I(N__20295));
    LocalMux I__2175 (
            .O(N__20301),
            .I(N__20290));
    Span4Mux_v I__2174 (
            .O(N__20298),
            .I(N__20290));
    LocalMux I__2173 (
            .O(N__20295),
            .I(pwm_duty_input_4));
    Odrv4 I__2172 (
            .O(N__20290),
            .I(pwm_duty_input_4));
    CascadeMux I__2171 (
            .O(N__20285),
            .I(N__20282));
    InMux I__2170 (
            .O(N__20282),
            .I(N__20278));
    InMux I__2169 (
            .O(N__20281),
            .I(N__20274));
    LocalMux I__2168 (
            .O(N__20278),
            .I(N__20271));
    InMux I__2167 (
            .O(N__20277),
            .I(N__20268));
    LocalMux I__2166 (
            .O(N__20274),
            .I(N__20265));
    Odrv4 I__2165 (
            .O(N__20271),
            .I(pwm_duty_input_5));
    LocalMux I__2164 (
            .O(N__20268),
            .I(pwm_duty_input_5));
    Odrv4 I__2163 (
            .O(N__20265),
            .I(pwm_duty_input_5));
    InMux I__2162 (
            .O(N__20258),
            .I(N__20255));
    LocalMux I__2161 (
            .O(N__20255),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ));
    InMux I__2160 (
            .O(N__20252),
            .I(N__20248));
    InMux I__2159 (
            .O(N__20251),
            .I(N__20245));
    LocalMux I__2158 (
            .O(N__20248),
            .I(N__20242));
    LocalMux I__2157 (
            .O(N__20245),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    Odrv4 I__2156 (
            .O(N__20242),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2155 (
            .O(N__20237),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    CascadeMux I__2154 (
            .O(N__20234),
            .I(N__20230));
    InMux I__2153 (
            .O(N__20233),
            .I(N__20225));
    InMux I__2152 (
            .O(N__20230),
            .I(N__20225));
    LocalMux I__2151 (
            .O(N__20225),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2150 (
            .O(N__20222),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2149 (
            .O(N__20219),
            .I(N__20213));
    InMux I__2148 (
            .O(N__20218),
            .I(N__20213));
    LocalMux I__2147 (
            .O(N__20213),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2146 (
            .O(N__20210),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    InMux I__2145 (
            .O(N__20207),
            .I(N__20201));
    InMux I__2144 (
            .O(N__20206),
            .I(N__20201));
    LocalMux I__2143 (
            .O(N__20201),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2142 (
            .O(N__20198),
            .I(bfn_3_20_0_));
    InMux I__2141 (
            .O(N__20195),
            .I(N__20189));
    InMux I__2140 (
            .O(N__20194),
            .I(N__20189));
    LocalMux I__2139 (
            .O(N__20189),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2138 (
            .O(N__20186),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2137 (
            .O(N__20183),
            .I(N__20177));
    InMux I__2136 (
            .O(N__20182),
            .I(N__20177));
    LocalMux I__2135 (
            .O(N__20177),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2134 (
            .O(N__20174),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2133 (
            .O(N__20171),
            .I(N__20167));
    InMux I__2132 (
            .O(N__20170),
            .I(N__20164));
    LocalMux I__2131 (
            .O(N__20167),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__2130 (
            .O(N__20164),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2129 (
            .O(N__20159),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2128 (
            .O(N__20156),
            .I(N__20150));
    InMux I__2127 (
            .O(N__20155),
            .I(N__20150));
    LocalMux I__2126 (
            .O(N__20150),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2125 (
            .O(N__20147),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2124 (
            .O(N__20144),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__2123 (
            .O(N__20141),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__2122 (
            .O(N__20138),
            .I(N__20134));
    InMux I__2121 (
            .O(N__20137),
            .I(N__20131));
    LocalMux I__2120 (
            .O(N__20134),
            .I(N__20128));
    LocalMux I__2119 (
            .O(N__20131),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    Odrv4 I__2118 (
            .O(N__20128),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2117 (
            .O(N__20123),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    CascadeMux I__2116 (
            .O(N__20120),
            .I(N__20117));
    InMux I__2115 (
            .O(N__20117),
            .I(N__20113));
    CascadeMux I__2114 (
            .O(N__20116),
            .I(N__20110));
    LocalMux I__2113 (
            .O(N__20113),
            .I(N__20107));
    InMux I__2112 (
            .O(N__20110),
            .I(N__20104));
    Odrv4 I__2111 (
            .O(N__20107),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    LocalMux I__2110 (
            .O(N__20104),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2109 (
            .O(N__20099),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    InMux I__2108 (
            .O(N__20096),
            .I(N__20090));
    InMux I__2107 (
            .O(N__20095),
            .I(N__20090));
    LocalMux I__2106 (
            .O(N__20090),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2105 (
            .O(N__20087),
            .I(bfn_3_19_0_));
    InMux I__2104 (
            .O(N__20084),
            .I(N__20078));
    InMux I__2103 (
            .O(N__20083),
            .I(N__20078));
    LocalMux I__2102 (
            .O(N__20078),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2101 (
            .O(N__20075),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2100 (
            .O(N__20072),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2099 (
            .O(N__20069),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__2098 (
            .O(N__20066),
            .I(N__20062));
    InMux I__2097 (
            .O(N__20065),
            .I(N__20059));
    LocalMux I__2096 (
            .O(N__20062),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    LocalMux I__2095 (
            .O(N__20059),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2094 (
            .O(N__20054),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__2093 (
            .O(N__20051),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2092 (
            .O(N__20048),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__2091 (
            .O(N__20045),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__2090 (
            .O(N__20042),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2089 (
            .O(N__20039),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    InMux I__2088 (
            .O(N__20036),
            .I(bfn_3_18_0_));
    InMux I__2087 (
            .O(N__20033),
            .I(N__20027));
    InMux I__2086 (
            .O(N__20032),
            .I(N__20027));
    LocalMux I__2085 (
            .O(N__20027),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2084 (
            .O(N__20024),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2083 (
            .O(N__20021),
            .I(N__20018));
    LocalMux I__2082 (
            .O(N__20018),
            .I(N__20014));
    InMux I__2081 (
            .O(N__20017),
            .I(N__20011));
    Odrv4 I__2080 (
            .O(N__20014),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    LocalMux I__2079 (
            .O(N__20011),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2078 (
            .O(N__20006),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    CascadeMux I__2077 (
            .O(N__20003),
            .I(N__20000));
    InMux I__2076 (
            .O(N__20000),
            .I(N__19997));
    LocalMux I__2075 (
            .O(N__19997),
            .I(N__19993));
    InMux I__2074 (
            .O(N__19996),
            .I(N__19990));
    Odrv4 I__2073 (
            .O(N__19993),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    LocalMux I__2072 (
            .O(N__19990),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2071 (
            .O(N__19985),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2070 (
            .O(N__19982),
            .I(N__19979));
    LocalMux I__2069 (
            .O(N__19979),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    CascadeMux I__2068 (
            .O(N__19976),
            .I(N__19973));
    InMux I__2067 (
            .O(N__19973),
            .I(N__19970));
    LocalMux I__2066 (
            .O(N__19970),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__2065 (
            .O(N__19967),
            .I(N__19964));
    LocalMux I__2064 (
            .O(N__19964),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__2063 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__2062 (
            .O(N__19958),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    CascadeMux I__2061 (
            .O(N__19955),
            .I(N__19952));
    InMux I__2060 (
            .O(N__19952),
            .I(N__19949));
    LocalMux I__2059 (
            .O(N__19949),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    CascadeMux I__2058 (
            .O(N__19946),
            .I(N__19943));
    InMux I__2057 (
            .O(N__19943),
            .I(N__19940));
    LocalMux I__2056 (
            .O(N__19940),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__2055 (
            .O(N__19937),
            .I(N__19934));
    LocalMux I__2054 (
            .O(N__19934),
            .I(N__19931));
    Span4Mux_s3_h I__2053 (
            .O(N__19931),
            .I(N__19928));
    Span4Mux_v I__2052 (
            .O(N__19928),
            .I(N__19925));
    Odrv4 I__2051 (
            .O(N__19925),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2050 (
            .O(N__19922),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2049 (
            .O(N__19919),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    CascadeMux I__2048 (
            .O(N__19916),
            .I(N__19913));
    InMux I__2047 (
            .O(N__19913),
            .I(N__19910));
    LocalMux I__2046 (
            .O(N__19910),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    CascadeMux I__2045 (
            .O(N__19907),
            .I(N__19904));
    InMux I__2044 (
            .O(N__19904),
            .I(N__19901));
    LocalMux I__2043 (
            .O(N__19901),
            .I(N__19897));
    CascadeMux I__2042 (
            .O(N__19900),
            .I(N__19894));
    Span4Mux_v I__2041 (
            .O(N__19897),
            .I(N__19891));
    InMux I__2040 (
            .O(N__19894),
            .I(N__19888));
    Sp12to4 I__2039 (
            .O(N__19891),
            .I(N__19883));
    LocalMux I__2038 (
            .O(N__19888),
            .I(N__19883));
    Span12Mux_h I__2037 (
            .O(N__19883),
            .I(N__19880));
    Odrv12 I__2036 (
            .O(N__19880),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    CascadeMux I__2035 (
            .O(N__19877),
            .I(N__19874));
    InMux I__2034 (
            .O(N__19874),
            .I(N__19871));
    LocalMux I__2033 (
            .O(N__19871),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__2032 (
            .O(N__19868),
            .I(N__19865));
    InMux I__2031 (
            .O(N__19865),
            .I(N__19862));
    LocalMux I__2030 (
            .O(N__19862),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__2029 (
            .O(N__19859),
            .I(N__19856));
    LocalMux I__2028 (
            .O(N__19856),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    CascadeMux I__2027 (
            .O(N__19853),
            .I(N__19850));
    InMux I__2026 (
            .O(N__19850),
            .I(N__19847));
    LocalMux I__2025 (
            .O(N__19847),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__2024 (
            .O(N__19844),
            .I(N__19841));
    LocalMux I__2023 (
            .O(N__19841),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    CascadeMux I__2022 (
            .O(N__19838),
            .I(N__19835));
    InMux I__2021 (
            .O(N__19835),
            .I(N__19832));
    LocalMux I__2020 (
            .O(N__19832),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__2019 (
            .O(N__19829),
            .I(N__19826));
    LocalMux I__2018 (
            .O(N__19826),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    CascadeMux I__2017 (
            .O(N__19823),
            .I(N__19819));
    CascadeMux I__2016 (
            .O(N__19822),
            .I(N__19815));
    InMux I__2015 (
            .O(N__19819),
            .I(N__19810));
    InMux I__2014 (
            .O(N__19818),
            .I(N__19810));
    InMux I__2013 (
            .O(N__19815),
            .I(N__19804));
    LocalMux I__2012 (
            .O(N__19810),
            .I(N__19800));
    InMux I__2011 (
            .O(N__19809),
            .I(N__19791));
    InMux I__2010 (
            .O(N__19808),
            .I(N__19791));
    InMux I__2009 (
            .O(N__19807),
            .I(N__19791));
    LocalMux I__2008 (
            .O(N__19804),
            .I(N__19788));
    InMux I__2007 (
            .O(N__19803),
            .I(N__19785));
    Span4Mux_v I__2006 (
            .O(N__19800),
            .I(N__19782));
    InMux I__2005 (
            .O(N__19799),
            .I(N__19779));
    InMux I__2004 (
            .O(N__19798),
            .I(N__19776));
    LocalMux I__2003 (
            .O(N__19791),
            .I(N__19769));
    Span4Mux_v I__2002 (
            .O(N__19788),
            .I(N__19769));
    LocalMux I__2001 (
            .O(N__19785),
            .I(N__19769));
    Odrv4 I__2000 (
            .O(N__19782),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    LocalMux I__1999 (
            .O(N__19779),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    LocalMux I__1998 (
            .O(N__19776),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    Odrv4 I__1997 (
            .O(N__19769),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    CascadeMux I__1996 (
            .O(N__19760),
            .I(\current_shift_inst.PI_CTRL.N_96_cascade_ ));
    InMux I__1995 (
            .O(N__19757),
            .I(N__19753));
    InMux I__1994 (
            .O(N__19756),
            .I(N__19750));
    LocalMux I__1993 (
            .O(N__19753),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    LocalMux I__1992 (
            .O(N__19750),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ));
    CascadeMux I__1991 (
            .O(N__19745),
            .I(N__19741));
    CascadeMux I__1990 (
            .O(N__19744),
            .I(N__19738));
    InMux I__1989 (
            .O(N__19741),
            .I(N__19732));
    InMux I__1988 (
            .O(N__19738),
            .I(N__19732));
    CascadeMux I__1987 (
            .O(N__19737),
            .I(N__19729));
    LocalMux I__1986 (
            .O(N__19732),
            .I(N__19726));
    InMux I__1985 (
            .O(N__19729),
            .I(N__19723));
    Odrv4 I__1984 (
            .O(N__19726),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    LocalMux I__1983 (
            .O(N__19723),
            .I(\current_shift_inst.PI_CTRL.control_out_2_0_3 ));
    InMux I__1982 (
            .O(N__19718),
            .I(N__19715));
    LocalMux I__1981 (
            .O(N__19715),
            .I(N__19711));
    InMux I__1980 (
            .O(N__19714),
            .I(N__19708));
    Span4Mux_s1_h I__1979 (
            .O(N__19711),
            .I(N__19705));
    LocalMux I__1978 (
            .O(N__19708),
            .I(pwm_duty_input_0));
    Odrv4 I__1977 (
            .O(N__19705),
            .I(pwm_duty_input_0));
    InMux I__1976 (
            .O(N__19700),
            .I(N__19696));
    InMux I__1975 (
            .O(N__19699),
            .I(N__19693));
    LocalMux I__1974 (
            .O(N__19696),
            .I(N__19690));
    LocalMux I__1973 (
            .O(N__19693),
            .I(pwm_duty_input_1));
    Odrv4 I__1972 (
            .O(N__19690),
            .I(pwm_duty_input_1));
    InMux I__1971 (
            .O(N__19685),
            .I(N__19682));
    LocalMux I__1970 (
            .O(N__19682),
            .I(N__19678));
    InMux I__1969 (
            .O(N__19681),
            .I(N__19675));
    Span4Mux_s1_h I__1968 (
            .O(N__19678),
            .I(N__19672));
    LocalMux I__1967 (
            .O(N__19675),
            .I(pwm_duty_input_2));
    Odrv4 I__1966 (
            .O(N__19672),
            .I(pwm_duty_input_2));
    CascadeMux I__1965 (
            .O(N__19667),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__1964 (
            .O(N__19664),
            .I(N__19661));
    LocalMux I__1963 (
            .O(N__19661),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    CascadeMux I__1962 (
            .O(N__19658),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ));
    InMux I__1961 (
            .O(N__19655),
            .I(N__19650));
    InMux I__1960 (
            .O(N__19654),
            .I(N__19645));
    InMux I__1959 (
            .O(N__19653),
            .I(N__19645));
    LocalMux I__1958 (
            .O(N__19650),
            .I(N__19642));
    LocalMux I__1957 (
            .O(N__19645),
            .I(pwm_duty_input_9));
    Odrv4 I__1956 (
            .O(N__19642),
            .I(pwm_duty_input_9));
    InMux I__1955 (
            .O(N__19637),
            .I(N__19632));
    InMux I__1954 (
            .O(N__19636),
            .I(N__19627));
    InMux I__1953 (
            .O(N__19635),
            .I(N__19627));
    LocalMux I__1952 (
            .O(N__19632),
            .I(N__19624));
    LocalMux I__1951 (
            .O(N__19627),
            .I(pwm_duty_input_7));
    Odrv4 I__1950 (
            .O(N__19624),
            .I(pwm_duty_input_7));
    CascadeMux I__1949 (
            .O(N__19619),
            .I(N__19614));
    InMux I__1948 (
            .O(N__19618),
            .I(N__19611));
    InMux I__1947 (
            .O(N__19617),
            .I(N__19608));
    InMux I__1946 (
            .O(N__19614),
            .I(N__19605));
    LocalMux I__1945 (
            .O(N__19611),
            .I(N__19602));
    LocalMux I__1944 (
            .O(N__19608),
            .I(pwm_duty_input_6));
    LocalMux I__1943 (
            .O(N__19605),
            .I(pwm_duty_input_6));
    Odrv4 I__1942 (
            .O(N__19602),
            .I(pwm_duty_input_6));
    InMux I__1941 (
            .O(N__19595),
            .I(N__19590));
    InMux I__1940 (
            .O(N__19594),
            .I(N__19587));
    InMux I__1939 (
            .O(N__19593),
            .I(N__19584));
    LocalMux I__1938 (
            .O(N__19590),
            .I(pwm_duty_input_8));
    LocalMux I__1937 (
            .O(N__19587),
            .I(pwm_duty_input_8));
    LocalMux I__1936 (
            .O(N__19584),
            .I(pwm_duty_input_8));
    CascadeMux I__1935 (
            .O(N__19577),
            .I(N__19574));
    InMux I__1934 (
            .O(N__19574),
            .I(N__19571));
    LocalMux I__1933 (
            .O(N__19571),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    CascadeMux I__1932 (
            .O(N__19568),
            .I(N__19565));
    InMux I__1931 (
            .O(N__19565),
            .I(N__19562));
    LocalMux I__1930 (
            .O(N__19562),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    CascadeMux I__1929 (
            .O(N__19559),
            .I(N__19556));
    InMux I__1928 (
            .O(N__19556),
            .I(N__19553));
    LocalMux I__1927 (
            .O(N__19553),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__1926 (
            .O(N__19550),
            .I(N__19547));
    LocalMux I__1925 (
            .O(N__19547),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__1924 (
            .O(N__19544),
            .I(N__19541));
    LocalMux I__1923 (
            .O(N__19541),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ));
    CascadeMux I__1922 (
            .O(N__19538),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    InMux I__1921 (
            .O(N__19535),
            .I(N__19532));
    LocalMux I__1920 (
            .O(N__19532),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    CascadeMux I__1919 (
            .O(N__19529),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ));
    InMux I__1918 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__1917 (
            .O(N__19523),
            .I(N__19520));
    Odrv4 I__1916 (
            .O(N__19520),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    InMux I__1915 (
            .O(N__19517),
            .I(N__19514));
    LocalMux I__1914 (
            .O(N__19514),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__1913 (
            .O(N__19511),
            .I(N__19504));
    InMux I__1912 (
            .O(N__19510),
            .I(N__19504));
    InMux I__1911 (
            .O(N__19509),
            .I(N__19501));
    LocalMux I__1910 (
            .O(N__19504),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__1909 (
            .O(N__19501),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__1908 (
            .O(N__19496),
            .I(N__19491));
    InMux I__1907 (
            .O(N__19495),
            .I(N__19485));
    InMux I__1906 (
            .O(N__19494),
            .I(N__19482));
    InMux I__1905 (
            .O(N__19491),
            .I(N__19475));
    InMux I__1904 (
            .O(N__19490),
            .I(N__19475));
    InMux I__1903 (
            .O(N__19489),
            .I(N__19475));
    CascadeMux I__1902 (
            .O(N__19488),
            .I(N__19472));
    LocalMux I__1901 (
            .O(N__19485),
            .I(N__19465));
    LocalMux I__1900 (
            .O(N__19482),
            .I(N__19465));
    LocalMux I__1899 (
            .O(N__19475),
            .I(N__19465));
    InMux I__1898 (
            .O(N__19472),
            .I(N__19461));
    Span4Mux_v I__1897 (
            .O(N__19465),
            .I(N__19458));
    InMux I__1896 (
            .O(N__19464),
            .I(N__19455));
    LocalMux I__1895 (
            .O(N__19461),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    Odrv4 I__1894 (
            .O(N__19458),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    LocalMux I__1893 (
            .O(N__19455),
            .I(\current_shift_inst.PI_CTRL.N_159 ));
    InMux I__1892 (
            .O(N__19448),
            .I(N__19436));
    InMux I__1891 (
            .O(N__19447),
            .I(N__19436));
    InMux I__1890 (
            .O(N__19446),
            .I(N__19436));
    InMux I__1889 (
            .O(N__19445),
            .I(N__19436));
    LocalMux I__1888 (
            .O(N__19436),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    CascadeMux I__1887 (
            .O(N__19433),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__1886 (
            .O(N__19430),
            .I(N__19427));
    LocalMux I__1885 (
            .O(N__19427),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__1884 (
            .O(N__19424),
            .I(N__19421));
    LocalMux I__1883 (
            .O(N__19421),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    CascadeMux I__1882 (
            .O(N__19418),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ));
    InMux I__1881 (
            .O(N__19415),
            .I(N__19412));
    LocalMux I__1880 (
            .O(N__19412),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__1879 (
            .O(N__19409),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ));
    InMux I__1878 (
            .O(N__19406),
            .I(N__19403));
    LocalMux I__1877 (
            .O(N__19403),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    CascadeMux I__1876 (
            .O(N__19400),
            .I(N__19397));
    InMux I__1875 (
            .O(N__19397),
            .I(N__19394));
    LocalMux I__1874 (
            .O(N__19394),
            .I(N__19391));
    Span4Mux_v I__1873 (
            .O(N__19391),
            .I(N__19388));
    Odrv4 I__1872 (
            .O(N__19388),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__1871 (
            .O(N__19385),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    CascadeMux I__1870 (
            .O(N__19382),
            .I(N__19379));
    InMux I__1869 (
            .O(N__19379),
            .I(N__19376));
    LocalMux I__1868 (
            .O(N__19376),
            .I(N__19373));
    Span4Mux_v I__1867 (
            .O(N__19373),
            .I(N__19370));
    Odrv4 I__1866 (
            .O(N__19370),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__1865 (
            .O(N__19367),
            .I(N__19364));
    LocalMux I__1864 (
            .O(N__19364),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__1863 (
            .O(N__19361),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    CascadeMux I__1862 (
            .O(N__19358),
            .I(N__19355));
    InMux I__1861 (
            .O(N__19355),
            .I(N__19352));
    LocalMux I__1860 (
            .O(N__19352),
            .I(N__19349));
    Span4Mux_h I__1859 (
            .O(N__19349),
            .I(N__19346));
    Odrv4 I__1858 (
            .O(N__19346),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__1857 (
            .O(N__19343),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__1856 (
            .O(N__19340),
            .I(N__19337));
    InMux I__1855 (
            .O(N__19337),
            .I(N__19334));
    LocalMux I__1854 (
            .O(N__19334),
            .I(N__19331));
    Odrv4 I__1853 (
            .O(N__19331),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__1852 (
            .O(N__19328),
            .I(N__19325));
    LocalMux I__1851 (
            .O(N__19325),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__1850 (
            .O(N__19322),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__1849 (
            .O(N__19319),
            .I(N__19316));
    InMux I__1848 (
            .O(N__19316),
            .I(N__19313));
    LocalMux I__1847 (
            .O(N__19313),
            .I(N__19310));
    Odrv4 I__1846 (
            .O(N__19310),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__1845 (
            .O(N__19307),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__1844 (
            .O(N__19304),
            .I(N__19301));
    LocalMux I__1843 (
            .O(N__19301),
            .I(N__19298));
    Odrv4 I__1842 (
            .O(N__19298),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    CascadeMux I__1841 (
            .O(N__19295),
            .I(N__19292));
    InMux I__1840 (
            .O(N__19292),
            .I(N__19289));
    LocalMux I__1839 (
            .O(N__19289),
            .I(N__19286));
    Span4Mux_v I__1838 (
            .O(N__19286),
            .I(N__19283));
    Odrv4 I__1837 (
            .O(N__19283),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ));
    InMux I__1836 (
            .O(N__19280),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__1835 (
            .O(N__19277),
            .I(N__19274));
    LocalMux I__1834 (
            .O(N__19274),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__1833 (
            .O(N__19271),
            .I(N__19268));
    LocalMux I__1832 (
            .O(N__19268),
            .I(N__19265));
    Span4Mux_v I__1831 (
            .O(N__19265),
            .I(N__19262));
    Odrv4 I__1830 (
            .O(N__19262),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    CascadeMux I__1829 (
            .O(N__19259),
            .I(N__19256));
    InMux I__1828 (
            .O(N__19256),
            .I(N__19253));
    LocalMux I__1827 (
            .O(N__19253),
            .I(N__19250));
    Odrv4 I__1826 (
            .O(N__19250),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__1825 (
            .O(N__19247),
            .I(N__19244));
    LocalMux I__1824 (
            .O(N__19244),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__1823 (
            .O(N__19241),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__1822 (
            .O(N__19238),
            .I(N__19235));
    InMux I__1821 (
            .O(N__19235),
            .I(N__19232));
    LocalMux I__1820 (
            .O(N__19232),
            .I(N__19229));
    Odrv4 I__1819 (
            .O(N__19229),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__1818 (
            .O(N__19226),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    CascadeMux I__1817 (
            .O(N__19223),
            .I(N__19220));
    InMux I__1816 (
            .O(N__19220),
            .I(N__19217));
    LocalMux I__1815 (
            .O(N__19217),
            .I(N__19214));
    Odrv4 I__1814 (
            .O(N__19214),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__1813 (
            .O(N__19211),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__1812 (
            .O(N__19208),
            .I(N__19205));
    InMux I__1811 (
            .O(N__19205),
            .I(N__19202));
    LocalMux I__1810 (
            .O(N__19202),
            .I(N__19199));
    Span4Mux_v I__1809 (
            .O(N__19199),
            .I(N__19196));
    Odrv4 I__1808 (
            .O(N__19196),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__1807 (
            .O(N__19193),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__1806 (
            .O(N__19190),
            .I(N__19187));
    InMux I__1805 (
            .O(N__19187),
            .I(N__19184));
    LocalMux I__1804 (
            .O(N__19184),
            .I(N__19181));
    Span4Mux_v I__1803 (
            .O(N__19181),
            .I(N__19178));
    Odrv4 I__1802 (
            .O(N__19178),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__1801 (
            .O(N__19175),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    CascadeMux I__1800 (
            .O(N__19172),
            .I(N__19169));
    InMux I__1799 (
            .O(N__19169),
            .I(N__19166));
    LocalMux I__1798 (
            .O(N__19166),
            .I(N__19163));
    Span4Mux_h I__1797 (
            .O(N__19163),
            .I(N__19160));
    Odrv4 I__1796 (
            .O(N__19160),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__1795 (
            .O(N__19157),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__1794 (
            .O(N__19154),
            .I(N__19151));
    InMux I__1793 (
            .O(N__19151),
            .I(N__19148));
    LocalMux I__1792 (
            .O(N__19148),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__1791 (
            .O(N__19145),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    CascadeMux I__1790 (
            .O(N__19142),
            .I(N__19139));
    InMux I__1789 (
            .O(N__19139),
            .I(N__19136));
    LocalMux I__1788 (
            .O(N__19136),
            .I(N__19133));
    Span4Mux_h I__1787 (
            .O(N__19133),
            .I(N__19130));
    Odrv4 I__1786 (
            .O(N__19130),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__1785 (
            .O(N__19127),
            .I(bfn_2_16_0_));
    CascadeMux I__1784 (
            .O(N__19124),
            .I(N__19121));
    InMux I__1783 (
            .O(N__19121),
            .I(N__19118));
    LocalMux I__1782 (
            .O(N__19118),
            .I(N__19115));
    Span4Mux_v I__1781 (
            .O(N__19115),
            .I(N__19112));
    Span4Mux_v I__1780 (
            .O(N__19112),
            .I(N__19109));
    Odrv4 I__1779 (
            .O(N__19109),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__1778 (
            .O(N__19106),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__1777 (
            .O(N__19103),
            .I(N__19100));
    InMux I__1776 (
            .O(N__19100),
            .I(N__19097));
    LocalMux I__1775 (
            .O(N__19097),
            .I(N__19094));
    Span4Mux_v I__1774 (
            .O(N__19094),
            .I(N__19091));
    Span4Mux_v I__1773 (
            .O(N__19091),
            .I(N__19088));
    Odrv4 I__1772 (
            .O(N__19088),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__1771 (
            .O(N__19085),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    CascadeMux I__1770 (
            .O(N__19082),
            .I(N__19079));
    InMux I__1769 (
            .O(N__19079),
            .I(N__19076));
    LocalMux I__1768 (
            .O(N__19076),
            .I(N__19073));
    Span4Mux_v I__1767 (
            .O(N__19073),
            .I(N__19070));
    Span4Mux_v I__1766 (
            .O(N__19070),
            .I(N__19067));
    Odrv4 I__1765 (
            .O(N__19067),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    CascadeMux I__1764 (
            .O(N__19064),
            .I(N__19061));
    InMux I__1763 (
            .O(N__19061),
            .I(N__19058));
    LocalMux I__1762 (
            .O(N__19058),
            .I(N__19055));
    Span4Mux_v I__1761 (
            .O(N__19055),
            .I(N__19052));
    Odrv4 I__1760 (
            .O(N__19052),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    InMux I__1759 (
            .O(N__19049),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__1758 (
            .O(N__19046),
            .I(N__19043));
    InMux I__1757 (
            .O(N__19043),
            .I(N__19040));
    LocalMux I__1756 (
            .O(N__19040),
            .I(N__19037));
    Span4Mux_v I__1755 (
            .O(N__19037),
            .I(N__19034));
    Span4Mux_v I__1754 (
            .O(N__19034),
            .I(N__19031));
    Odrv4 I__1753 (
            .O(N__19031),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__1752 (
            .O(N__19028),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    CascadeMux I__1751 (
            .O(N__19025),
            .I(N__19022));
    InMux I__1750 (
            .O(N__19022),
            .I(N__19019));
    LocalMux I__1749 (
            .O(N__19019),
            .I(N__19016));
    Span4Mux_v I__1748 (
            .O(N__19016),
            .I(N__19013));
    Span4Mux_v I__1747 (
            .O(N__19013),
            .I(N__19010));
    Odrv4 I__1746 (
            .O(N__19010),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__1745 (
            .O(N__19007),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__1744 (
            .O(N__19004),
            .I(N__19001));
    InMux I__1743 (
            .O(N__19001),
            .I(N__18998));
    LocalMux I__1742 (
            .O(N__18998),
            .I(N__18995));
    Span4Mux_v I__1741 (
            .O(N__18995),
            .I(N__18992));
    Span4Mux_v I__1740 (
            .O(N__18992),
            .I(N__18989));
    Odrv4 I__1739 (
            .O(N__18989),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__1738 (
            .O(N__18986),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__1737 (
            .O(N__18983),
            .I(N__18980));
    InMux I__1736 (
            .O(N__18980),
            .I(N__18977));
    LocalMux I__1735 (
            .O(N__18977),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__1734 (
            .O(N__18974),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    CascadeMux I__1733 (
            .O(N__18971),
            .I(N__18968));
    InMux I__1732 (
            .O(N__18968),
            .I(N__18965));
    LocalMux I__1731 (
            .O(N__18965),
            .I(N__18962));
    Span4Mux_h I__1730 (
            .O(N__18962),
            .I(N__18959));
    Odrv4 I__1729 (
            .O(N__18959),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__1728 (
            .O(N__18956),
            .I(bfn_2_15_0_));
    CascadeMux I__1727 (
            .O(N__18953),
            .I(N__18950));
    InMux I__1726 (
            .O(N__18950),
            .I(N__18947));
    LocalMux I__1725 (
            .O(N__18947),
            .I(N__18944));
    Span4Mux_v I__1724 (
            .O(N__18944),
            .I(N__18941));
    Span4Mux_v I__1723 (
            .O(N__18941),
            .I(N__18938));
    Odrv4 I__1722 (
            .O(N__18938),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__1721 (
            .O(N__18935),
            .I(N__18932));
    LocalMux I__1720 (
            .O(N__18932),
            .I(N__18929));
    Span4Mux_v I__1719 (
            .O(N__18929),
            .I(N__18926));
    Odrv4 I__1718 (
            .O(N__18926),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__1717 (
            .O(N__18923),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    CascadeMux I__1716 (
            .O(N__18920),
            .I(N__18917));
    InMux I__1715 (
            .O(N__18917),
            .I(N__18914));
    LocalMux I__1714 (
            .O(N__18914),
            .I(N__18911));
    Span4Mux_s3_h I__1713 (
            .O(N__18911),
            .I(N__18908));
    Span4Mux_v I__1712 (
            .O(N__18908),
            .I(N__18905));
    Span4Mux_v I__1711 (
            .O(N__18905),
            .I(N__18902));
    Odrv4 I__1710 (
            .O(N__18902),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__1709 (
            .O(N__18899),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__1708 (
            .O(N__18896),
            .I(N__18893));
    InMux I__1707 (
            .O(N__18893),
            .I(N__18890));
    LocalMux I__1706 (
            .O(N__18890),
            .I(N__18887));
    Span4Mux_v I__1705 (
            .O(N__18887),
            .I(N__18884));
    Span4Mux_v I__1704 (
            .O(N__18884),
            .I(N__18881));
    Odrv4 I__1703 (
            .O(N__18881),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    CascadeMux I__1702 (
            .O(N__18878),
            .I(N__18875));
    InMux I__1701 (
            .O(N__18875),
            .I(N__18872));
    LocalMux I__1700 (
            .O(N__18872),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__1699 (
            .O(N__18869),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    CascadeMux I__1698 (
            .O(N__18866),
            .I(N__18863));
    InMux I__1697 (
            .O(N__18863),
            .I(N__18860));
    LocalMux I__1696 (
            .O(N__18860),
            .I(N__18857));
    Span4Mux_v I__1695 (
            .O(N__18857),
            .I(N__18854));
    Span4Mux_v I__1694 (
            .O(N__18854),
            .I(N__18851));
    Odrv4 I__1693 (
            .O(N__18851),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__1692 (
            .O(N__18848),
            .I(N__18845));
    LocalMux I__1691 (
            .O(N__18845),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__1690 (
            .O(N__18842),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__1689 (
            .O(N__18839),
            .I(N__18836));
    InMux I__1688 (
            .O(N__18836),
            .I(N__18833));
    LocalMux I__1687 (
            .O(N__18833),
            .I(N__18830));
    Span4Mux_v I__1686 (
            .O(N__18830),
            .I(N__18827));
    Span4Mux_v I__1685 (
            .O(N__18827),
            .I(N__18824));
    Odrv4 I__1684 (
            .O(N__18824),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__1683 (
            .O(N__18821),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__1682 (
            .O(N__18818),
            .I(N__18815));
    InMux I__1681 (
            .O(N__18815),
            .I(N__18812));
    LocalMux I__1680 (
            .O(N__18812),
            .I(N__18809));
    Span12Mux_v I__1679 (
            .O(N__18809),
            .I(N__18806));
    Odrv12 I__1678 (
            .O(N__18806),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__1677 (
            .O(N__18803),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__1676 (
            .O(N__18800),
            .I(N__18797));
    InMux I__1675 (
            .O(N__18797),
            .I(N__18794));
    LocalMux I__1674 (
            .O(N__18794),
            .I(N__18791));
    Span4Mux_v I__1673 (
            .O(N__18791),
            .I(N__18788));
    Span4Mux_v I__1672 (
            .O(N__18788),
            .I(N__18785));
    Odrv4 I__1671 (
            .O(N__18785),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__1670 (
            .O(N__18782),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    CascadeMux I__1669 (
            .O(N__18779),
            .I(N__18776));
    InMux I__1668 (
            .O(N__18776),
            .I(N__18773));
    LocalMux I__1667 (
            .O(N__18773),
            .I(N__18770));
    Span12Mux_h I__1666 (
            .O(N__18770),
            .I(N__18767));
    Odrv12 I__1665 (
            .O(N__18767),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    InMux I__1664 (
            .O(N__18764),
            .I(bfn_2_14_0_));
    InMux I__1663 (
            .O(N__18761),
            .I(N__18758));
    LocalMux I__1662 (
            .O(N__18758),
            .I(N__18755));
    Odrv4 I__1661 (
            .O(N__18755),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    InMux I__1660 (
            .O(N__18752),
            .I(N__18749));
    LocalMux I__1659 (
            .O(N__18749),
            .I(N_42_i_i));
    InMux I__1658 (
            .O(N__18746),
            .I(N__18743));
    LocalMux I__1657 (
            .O(N__18743),
            .I(un7_start_stop_0_a2));
    InMux I__1656 (
            .O(N__18740),
            .I(N__18737));
    LocalMux I__1655 (
            .O(N__18737),
            .I(N__18734));
    Odrv4 I__1654 (
            .O(N__18734),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    InMux I__1653 (
            .O(N__18731),
            .I(N__18722));
    InMux I__1652 (
            .O(N__18730),
            .I(N__18722));
    InMux I__1651 (
            .O(N__18729),
            .I(N__18722));
    LocalMux I__1650 (
            .O(N__18722),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__1649 (
            .O(N__18719),
            .I(N__18716));
    LocalMux I__1648 (
            .O(N__18716),
            .I(N__18713));
    Odrv4 I__1647 (
            .O(N__18713),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__1646 (
            .O(N__18710),
            .I(N__18707));
    LocalMux I__1645 (
            .O(N__18707),
            .I(N__18704));
    Odrv4 I__1644 (
            .O(N__18704),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__1643 (
            .O(N__18701),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__1642 (
            .O(N__18698),
            .I(N__18695));
    LocalMux I__1641 (
            .O(N__18695),
            .I(N__18692));
    Odrv4 I__1640 (
            .O(N__18692),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    InMux I__1639 (
            .O(N__18689),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__1638 (
            .O(N__18686),
            .I(N__18683));
    LocalMux I__1637 (
            .O(N__18683),
            .I(N__18680));
    Odrv4 I__1636 (
            .O(N__18680),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    InMux I__1635 (
            .O(N__18677),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    InMux I__1634 (
            .O(N__18674),
            .I(N__18671));
    LocalMux I__1633 (
            .O(N__18671),
            .I(N__18668));
    Span4Mux_h I__1632 (
            .O(N__18668),
            .I(N__18665));
    Odrv4 I__1631 (
            .O(N__18665),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    CascadeMux I__1630 (
            .O(N__18662),
            .I(N__18649));
    CascadeMux I__1629 (
            .O(N__18661),
            .I(N__18646));
    CascadeMux I__1628 (
            .O(N__18660),
            .I(N__18643));
    CascadeMux I__1627 (
            .O(N__18659),
            .I(N__18640));
    CascadeMux I__1626 (
            .O(N__18658),
            .I(N__18637));
    CascadeMux I__1625 (
            .O(N__18657),
            .I(N__18634));
    CascadeMux I__1624 (
            .O(N__18656),
            .I(N__18631));
    CascadeMux I__1623 (
            .O(N__18655),
            .I(N__18628));
    CascadeMux I__1622 (
            .O(N__18654),
            .I(N__18625));
    CascadeMux I__1621 (
            .O(N__18653),
            .I(N__18622));
    InMux I__1620 (
            .O(N__18652),
            .I(N__18618));
    InMux I__1619 (
            .O(N__18649),
            .I(N__18609));
    InMux I__1618 (
            .O(N__18646),
            .I(N__18609));
    InMux I__1617 (
            .O(N__18643),
            .I(N__18609));
    InMux I__1616 (
            .O(N__18640),
            .I(N__18609));
    InMux I__1615 (
            .O(N__18637),
            .I(N__18606));
    InMux I__1614 (
            .O(N__18634),
            .I(N__18599));
    InMux I__1613 (
            .O(N__18631),
            .I(N__18599));
    InMux I__1612 (
            .O(N__18628),
            .I(N__18599));
    InMux I__1611 (
            .O(N__18625),
            .I(N__18592));
    InMux I__1610 (
            .O(N__18622),
            .I(N__18592));
    InMux I__1609 (
            .O(N__18621),
            .I(N__18592));
    LocalMux I__1608 (
            .O(N__18618),
            .I(N__18585));
    LocalMux I__1607 (
            .O(N__18609),
            .I(N__18585));
    LocalMux I__1606 (
            .O(N__18606),
            .I(N__18585));
    LocalMux I__1605 (
            .O(N__18599),
            .I(N__18580));
    LocalMux I__1604 (
            .O(N__18592),
            .I(N__18580));
    Span4Mux_v I__1603 (
            .O(N__18585),
            .I(N__18575));
    Span4Mux_v I__1602 (
            .O(N__18580),
            .I(N__18575));
    Odrv4 I__1601 (
            .O(N__18575),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    InMux I__1600 (
            .O(N__18572),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__1599 (
            .O(N__18569),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    InMux I__1598 (
            .O(N__18566),
            .I(N__18563));
    LocalMux I__1597 (
            .O(N__18563),
            .I(N__18560));
    Span4Mux_v I__1596 (
            .O(N__18560),
            .I(N__18557));
    Odrv4 I__1595 (
            .O(N__18557),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__1594 (
            .O(N__18554),
            .I(N__18551));
    InMux I__1593 (
            .O(N__18551),
            .I(N__18548));
    LocalMux I__1592 (
            .O(N__18548),
            .I(N__18545));
    Span4Mux_v I__1591 (
            .O(N__18545),
            .I(N__18542));
    Span4Mux_v I__1590 (
            .O(N__18542),
            .I(N__18539));
    Odrv4 I__1589 (
            .O(N__18539),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__1588 (
            .O(N__18536),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    CascadeMux I__1587 (
            .O(N__18533),
            .I(N__18530));
    InMux I__1586 (
            .O(N__18530),
            .I(N__18527));
    LocalMux I__1585 (
            .O(N__18527),
            .I(N__18524));
    Odrv4 I__1584 (
            .O(N__18524),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    InMux I__1583 (
            .O(N__18521),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    InMux I__1582 (
            .O(N__18518),
            .I(N__18515));
    LocalMux I__1581 (
            .O(N__18515),
            .I(N__18512));
    Odrv4 I__1580 (
            .O(N__18512),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    InMux I__1579 (
            .O(N__18509),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__1578 (
            .O(N__18506),
            .I(N__18503));
    LocalMux I__1577 (
            .O(N__18503),
            .I(N__18500));
    Odrv4 I__1576 (
            .O(N__18500),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    InMux I__1575 (
            .O(N__18497),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    InMux I__1574 (
            .O(N__18494),
            .I(N__18491));
    LocalMux I__1573 (
            .O(N__18491),
            .I(N__18488));
    Odrv4 I__1572 (
            .O(N__18488),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__1571 (
            .O(N__18485),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    InMux I__1570 (
            .O(N__18482),
            .I(N__18479));
    LocalMux I__1569 (
            .O(N__18479),
            .I(N__18476));
    Span4Mux_v I__1568 (
            .O(N__18476),
            .I(N__18473));
    Odrv4 I__1567 (
            .O(N__18473),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    InMux I__1566 (
            .O(N__18470),
            .I(bfn_1_14_0_));
    InMux I__1565 (
            .O(N__18467),
            .I(N__18464));
    LocalMux I__1564 (
            .O(N__18464),
            .I(N__18461));
    Span4Mux_v I__1563 (
            .O(N__18461),
            .I(N__18458));
    Odrv4 I__1562 (
            .O(N__18458),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    InMux I__1561 (
            .O(N__18455),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    InMux I__1560 (
            .O(N__18452),
            .I(N__18449));
    LocalMux I__1559 (
            .O(N__18449),
            .I(N__18446));
    Odrv4 I__1558 (
            .O(N__18446),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__1557 (
            .O(N__18443),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__1556 (
            .O(N__18440),
            .I(N__18437));
    LocalMux I__1555 (
            .O(N__18437),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    InMux I__1554 (
            .O(N__18434),
            .I(N__18431));
    LocalMux I__1553 (
            .O(N__18431),
            .I(N__18428));
    Span4Mux_v I__1552 (
            .O(N__18428),
            .I(N__18425));
    Odrv4 I__1551 (
            .O(N__18425),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__1550 (
            .O(N__18422),
            .I(N__18419));
    InMux I__1549 (
            .O(N__18419),
            .I(N__18416));
    LocalMux I__1548 (
            .O(N__18416),
            .I(N__18413));
    Span4Mux_v I__1547 (
            .O(N__18413),
            .I(N__18410));
    Odrv4 I__1546 (
            .O(N__18410),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    InMux I__1545 (
            .O(N__18407),
            .I(N__18404));
    LocalMux I__1544 (
            .O(N__18404),
            .I(N__18401));
    Span4Mux_v I__1543 (
            .O(N__18401),
            .I(N__18398));
    Odrv4 I__1542 (
            .O(N__18398),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__1541 (
            .O(N__18395),
            .I(N__18392));
    InMux I__1540 (
            .O(N__18392),
            .I(N__18389));
    LocalMux I__1539 (
            .O(N__18389),
            .I(N__18386));
    Span4Mux_v I__1538 (
            .O(N__18386),
            .I(N__18383));
    Odrv4 I__1537 (
            .O(N__18383),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    InMux I__1536 (
            .O(N__18380),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__1535 (
            .O(N__18377),
            .I(N__18374));
    LocalMux I__1534 (
            .O(N__18374),
            .I(N__18371));
    Span4Mux_h I__1533 (
            .O(N__18371),
            .I(N__18368));
    Odrv4 I__1532 (
            .O(N__18368),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__1531 (
            .O(N__18365),
            .I(N__18362));
    InMux I__1530 (
            .O(N__18362),
            .I(N__18359));
    LocalMux I__1529 (
            .O(N__18359),
            .I(N__18356));
    Span4Mux_v I__1528 (
            .O(N__18356),
            .I(N__18353));
    Odrv4 I__1527 (
            .O(N__18353),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    InMux I__1526 (
            .O(N__18350),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    IoInMux I__1525 (
            .O(N__18347),
            .I(N__18344));
    LocalMux I__1524 (
            .O(N__18344),
            .I(N__18341));
    Span4Mux_s3_v I__1523 (
            .O(N__18341),
            .I(N__18338));
    Span4Mux_h I__1522 (
            .O(N__18338),
            .I(N__18335));
    Sp12to4 I__1521 (
            .O(N__18335),
            .I(N__18332));
    Span12Mux_v I__1520 (
            .O(N__18332),
            .I(N__18329));
    Span12Mux_v I__1519 (
            .O(N__18329),
            .I(N__18326));
    Odrv12 I__1518 (
            .O(N__18326),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1517 (
            .O(N__18323),
            .I(N__18320));
    LocalMux I__1516 (
            .O(N__18320),
            .I(N__18317));
    IoSpan4Mux I__1515 (
            .O(N__18317),
            .I(N__18314));
    IoSpan4Mux I__1514 (
            .O(N__18314),
            .I(N__18311));
    Odrv4 I__1513 (
            .O(N__18311),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_3_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_24_0_));
    defparam IN_MUX_bfv_3_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_25_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_3_25_0_));
    defparam IN_MUX_bfv_3_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_26_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_3_26_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_3_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_3_20_0_));
    defparam IN_MUX_bfv_4_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_23_0_));
    defparam IN_MUX_bfv_4_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_24_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_4_24_0_));
    defparam IN_MUX_bfv_4_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_25_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_4_25_0_));
    defparam IN_MUX_bfv_7_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_23_0_));
    defparam IN_MUX_bfv_7_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_24_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_7_24_0_));
    defparam IN_MUX_bfv_5_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_25_0_));
    defparam IN_MUX_bfv_5_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_26_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_5_26_0_));
    defparam IN_MUX_bfv_5_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_27_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_5_27_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_10_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_24_0_));
    defparam IN_MUX_bfv_10_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_25_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_10_25_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_10_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_7_0_));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_10_8_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_12_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_12_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_10_13_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_15_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_15_21_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_8_20_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18347),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__18323),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__33686),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_162_i_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0  (
            .USERSIGNALTOGLOBALBUFFER(N__34180),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un1_start_g ));
    ICE_GB \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0  (
            .USERSIGNALTOGLOBALBUFFER(N__32198),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_hc.un1_start_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__38001),
            .CLKHFEN(N__38003),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__38002),
            .RGB2PWM(N__18752),
            .RGB1(rgb_g),
            .CURREN(N__37975),
            .RGB2(rgb_b),
            .RGB1PWM(N__18746),
            .RGB0PWM(N__46961),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__18440),
            .in2(_gnd_net_),
            .in3(N__18652),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__18434),
            .in2(N__18422),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__18407),
            .in2(N__18395),
            .in3(N__18380),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__18377),
            .in2(N__18365),
            .in3(N__18350),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__18566),
            .in2(N__18554),
            .in3(N__18536),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__18621),
            .in2(N__18533),
            .in3(N__18521),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__18518),
            .in2(N__18653),
            .in3(N__18509),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__18506),
            .in2(N__18658),
            .in3(N__18497),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__18494),
            .in2(N__18654),
            .in3(N__18485),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__18482),
            .in2(N__18659),
            .in3(N__18470),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__18467),
            .in2(N__18655),
            .in3(N__18455),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__18452),
            .in2(N__18660),
            .in3(N__18443),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__18710),
            .in2(N__18656),
            .in3(N__18701),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__18698),
            .in2(N__18661),
            .in3(N__18689),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__18686),
            .in2(N__18657),
            .in3(N__18677),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__18674),
            .in2(N__18662),
            .in3(N__18572),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18569),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_1_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_1_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_1_15_2 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_1_15_2  (
            .in0(N__23064),
            .in1(N__23255),
            .in2(N__22634),
            .in3(N__19328),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47673),
            .ce(),
            .sr(N__46919));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_1_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_1_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_1_15_4 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_1_15_4  (
            .in0(N__23063),
            .in1(N__23254),
            .in2(N__22633),
            .in3(N__19247),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47673),
            .ce(),
            .sr(N__46919));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_1_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_1_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_1_16_3 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_1_16_3  (
            .in0(N__23181),
            .in1(N__23077),
            .in2(N__19064),
            .in3(N__22598),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47662),
            .ce(),
            .sr(N__46923));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_6 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_6  (
            .in0(N__22597),
            .in1(N__23182),
            .in2(N__23084),
            .in3(N__19367),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47662),
            .ce(),
            .sr(N__46923));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_1_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_1_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_1_17_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_1_17_1  (
            .in0(N__18935),
            .in1(N__23076),
            .in2(_gnd_net_),
            .in3(N__22609),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47652),
            .ce(),
            .sr(N__46927));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_1_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_1_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_1_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24997),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47639),
            .ce(),
            .sr(N__46931));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18740),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47617),
            .ce(),
            .sr(N__46936));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_1_21_0  (
            .in0(N__19511),
            .in1(N__43843),
            .in2(_gnd_net_),
            .in3(N__19799),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_5 .LUT_INIT=16'b0100010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_21_5  (
            .in0(N__43844),
            .in1(N__19798),
            .in2(N__20686),
            .in3(N__19510),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2  (
            .in0(N__19818),
            .in1(N__43845),
            .in2(N__19488),
            .in3(N__20462),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47596),
            .ce(),
            .sr(N__46937));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_22_3  (
            .in0(N__18731),
            .in1(N__19937),
            .in2(N__19745),
            .in3(N__19448),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47596),
            .ce(),
            .sr(N__46937));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_22_4  (
            .in0(N__19445),
            .in1(N__19271),
            .in2(N__19737),
            .in3(N__18730),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47596),
            .ce(),
            .sr(N__46937));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_5 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_22_5  (
            .in0(N__18729),
            .in1(N__18719),
            .in2(N__19744),
            .in3(N__19447),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47596),
            .ce(),
            .sr(N__46937));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_6 .LUT_INIT=16'b1101110011011101;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_6  (
            .in0(N__19446),
            .in1(N__20645),
            .in2(N__19823),
            .in3(N__19757),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47596),
            .ce(),
            .sr(N__46937));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_0 .LUT_INIT=16'b1100111100001010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_23_0  (
            .in0(N__19807),
            .in1(N__19490),
            .in2(N__43855),
            .in3(N__20393),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47589),
            .ce(),
            .sr(N__46939));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_23_1 .LUT_INIT=16'b1010000011111100;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_23_1  (
            .in0(N__19489),
            .in1(N__19808),
            .in2(N__20498),
            .in3(N__43846),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47589),
            .ce(),
            .sr(N__46939));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_23_3 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_23_3  (
            .in0(N__20687),
            .in1(N__18761),
            .in2(N__20363),
            .in3(N__19495),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47589),
            .ce(),
            .sr(N__46939));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_5 .LUT_INIT=16'b1010000011101110;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_23_5  (
            .in0(N__20429),
            .in1(N__19809),
            .in2(N__19496),
            .in3(N__43847),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47589),
            .ce(),
            .sr(N__46939));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_24_1 .LUT_INIT=16'b1000100011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_24_1  (
            .in0(N__20525),
            .in1(N__19494),
            .in2(N__19822),
            .in3(N__43851),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47583),
            .ce(),
            .sr(N__46940));
    defparam \phase_controller_inst1.N_42_i_i_LC_1_30_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.N_42_i_i_LC_1_30_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.N_42_i_i_LC_1_30_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \phase_controller_inst1.N_42_i_i_LC_1_30_5  (
            .in0(N__30826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46959),
            .lcout(N_42_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.un7_start_stop_0_a2_LC_1_30_6  (
            .in0(N__46960),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30827),
            .lcout(un7_start_stop_0_a2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_2_12_5 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_2_12_5  (
            .in0(N__23082),
            .in1(N__23223),
            .in2(N__18878),
            .in3(N__22602),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47694),
            .ce(),
            .sr(N__46903));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_2_12_6 .LUT_INIT=16'b1100010011000101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_2_12_6  (
            .in0(N__23222),
            .in1(N__18848),
            .in2(N__22631),
            .in3(N__23083),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47694),
            .ce(),
            .sr(N__46903));
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__20824),
            .in2(N__19900),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__20880),
            .in2(N__18953),
            .in3(N__18923),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__22862),
            .in2(N__18920),
            .in3(N__18899),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__22766),
            .in2(N__18896),
            .in3(N__18869),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__22820),
            .in2(N__18866),
            .in3(N__18842),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__20787),
            .in2(N__18839),
            .in3(N__18821),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__22912),
            .in2(N__18818),
            .in3(N__18803),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__21244),
            .in2(N__18800),
            .in3(N__18782),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__23287),
            .in2(N__18779),
            .in3(N__18764),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__21119),
            .in2(N__19124),
            .in3(N__19106),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__21356),
            .in2(N__19103),
            .in3(N__19085),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__21296),
            .in2(N__19082),
            .in3(N__19049),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__21157),
            .in2(N__19046),
            .in3(N__19028),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_2_14_5  (
            .in0(_gnd_net_),
            .in1(N__21389),
            .in2(N__19025),
            .in3(N__19007),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__21187),
            .in2(N__19004),
            .in3(N__18986),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__21090),
            .in2(N__18983),
            .in3(N__18974),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__20974),
            .in2(N__18971),
            .in3(N__18956),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__21032),
            .in2(N__19259),
            .in3(N__19241),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__21061),
            .in2(N__19238),
            .in3(N__19226),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__21570),
            .in2(N__19223),
            .in3(N__19211),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__20947),
            .in2(N__19208),
            .in3(N__19193),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__21005),
            .in2(N__19190),
            .in3(N__19175),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__22695),
            .in2(N__19172),
            .in3(N__19157),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__21597),
            .in2(N__19154),
            .in3(N__19145),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__21462),
            .in2(N__19142),
            .in3(N__19127),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__21517),
            .in2(N__19400),
            .in3(N__19385),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__21423),
            .in2(N__19382),
            .in3(N__19361),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__21493),
            .in2(N__19358),
            .in3(N__19343),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__22727),
            .in2(N__19340),
            .in3(N__19322),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(N__21334),
            .in2(N__19319),
            .in3(N__19307),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_16_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_2_16_6  (
            .in0(N__19304),
            .in1(N__23159),
            .in2(N__19295),
            .in3(N__19280),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_2_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_2_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_2_17_1 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_2_17_1  (
            .in0(N__23081),
            .in1(N__23189),
            .in2(N__22632),
            .in3(N__19277),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47641),
            .ce(),
            .sr(N__46924));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_18_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_2_18_4  (
            .in0(_gnd_net_),
            .in1(N__21637),
            .in2(_gnd_net_),
            .in3(N__20845),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47628),
            .ce(),
            .sr(N__46928));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_19_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_19_0  (
            .in0(_gnd_net_),
            .in1(N__20379),
            .in2(_gnd_net_),
            .in3(N__20484),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_2  (
            .in0(N__20219),
            .in1(N__20581),
            .in2(N__20549),
            .in3(N__20233),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_3  (
            .in0(_gnd_net_),
            .in1(N__19996),
            .in2(_gnd_net_),
            .in3(N__20032),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_4  (
            .in0(N__20170),
            .in1(N__20017),
            .in2(N__19433),
            .in3(N__19430),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6  (
            .in0(N__20033),
            .in1(N__20156),
            .in2(N__20116),
            .in3(N__20137),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_7  (
            .in0(N__20155),
            .in1(N__20218),
            .in2(N__20234),
            .in3(N__20065),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_20_0  (
            .in0(N__20021),
            .in1(N__19424),
            .in2(N__20003),
            .in3(N__19550),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_2_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_2_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_2_20_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIQP82_27_LC_2_20_1  (
            .in0(_gnd_net_),
            .in1(N__20704),
            .in2(_gnd_net_),
            .in3(N__20183),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_9_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_2_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_2_20_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_21_LC_2_20_2  (
            .in0(N__20171),
            .in1(N__20251),
            .in2(N__19418),
            .in3(N__20066),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_3  (
            .in0(N__19415),
            .in1(N__19517),
            .in2(N__19409),
            .in3(N__19406),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_4  (
            .in0(_gnd_net_),
            .in1(N__20083),
            .in2(_gnd_net_),
            .in3(N__20095),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_5 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_0_6_LC_2_20_5  (
            .in0(N__20524),
            .in1(N__19544),
            .in2(N__20461),
            .in3(N__20418),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_6  (
            .in0(N__20182),
            .in1(N__20084),
            .in2(N__20705),
            .in3(N__20096),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_2_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_2_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_2_21_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_2_21_1  (
            .in0(N__20138),
            .in1(_gnd_net_),
            .in2(N__20120),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_2_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_2_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_2_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_2_21_2  (
            .in0(N__20194),
            .in1(N__20206),
            .in2(N__19538),
            .in3(N__20252),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_2_21_3  (
            .in0(N__19535),
            .in1(N__20531),
            .in2(N__19529),
            .in3(N__19526),
            .lcout(\current_shift_inst.PI_CTRL.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_21_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_21_5  (
            .in0(N__20207),
            .in1(N__20563),
            .in2(N__20606),
            .in3(N__20195),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_21_7 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISN3A1_4_LC_2_21_7  (
            .in0(N__20679),
            .in1(N__43804),
            .in2(_gnd_net_),
            .in3(N__19509),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_6 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_6  (
            .in0(N__19464),
            .in1(N__20612),
            .in2(N__20356),
            .in3(N__43821),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(\current_shift_inst.PI_CTRL.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_22_7 .LUT_INIT=16'b0101000101010000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI8OCG4_3_LC_2_22_7  (
            .in0(N__20641),
            .in1(N__19803),
            .in2(N__19760),
            .in3(N__19756),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_23_2  (
            .in0(N__19714),
            .in1(N__19699),
            .in2(_gnd_net_),
            .in3(N__19681),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_23_3  (
            .in0(_gnd_net_),
            .in1(N__19636),
            .in2(_gnd_net_),
            .in3(N__20277),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_23_4  (
            .in0(N__19617),
            .in1(N__19595),
            .in2(N__19667),
            .in3(N__19654),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_5 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_5  (
            .in0(N__19664),
            .in1(N__20328),
            .in2(N__19658),
            .in3(N__20304),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_7  (
            .in0(N__19653),
            .in1(N__19635),
            .in2(N__19619),
            .in3(N__19594),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_0 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_3_14_0  (
            .in0(N__23228),
            .in1(N__23047),
            .in2(N__19577),
            .in3(N__22629),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47663),
            .ce(),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_3_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_3_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_3_14_1 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_3_14_1  (
            .in0(N__22624),
            .in1(N__23230),
            .in2(N__19568),
            .in3(N__23051),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47663),
            .ce(),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_3 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_3_14_3  (
            .in0(N__22626),
            .in1(N__23232),
            .in2(N__19559),
            .in3(N__23053),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47663),
            .ce(),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_4 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_3_14_4  (
            .in0(N__23229),
            .in1(N__23048),
            .in2(N__19916),
            .in3(N__22630),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47663),
            .ce(),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5 .LUT_INIT=16'b0011110000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_3_14_5  (
            .in0(N__22627),
            .in1(N__20834),
            .in2(N__19907),
            .in3(N__23054),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47663),
            .ce(),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_3_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_3_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_3_14_6 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_3_14_6  (
            .in0(N__23227),
            .in1(N__23046),
            .in2(N__19877),
            .in3(N__22628),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47663),
            .ce(),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_3_14_7 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_3_14_7  (
            .in0(N__22625),
            .in1(N__23231),
            .in2(N__19868),
            .in3(N__23052),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47663),
            .ce(),
            .sr(N__46907));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_3_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_3_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_3_15_1 .LUT_INIT=16'b1101110011011000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_3_15_1  (
            .in0(N__22615),
            .in1(N__19859),
            .in2(N__23259),
            .in3(N__23039),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47653),
            .ce(),
            .sr(N__46911));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_4 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_3_15_4  (
            .in0(N__23035),
            .in1(N__23234),
            .in2(N__19853),
            .in3(N__22616),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47653),
            .ce(),
            .sr(N__46911));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_5 .LUT_INIT=16'b1101110011011000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_3_15_5  (
            .in0(N__22614),
            .in1(N__19844),
            .in2(N__23258),
            .in3(N__23038),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47653),
            .ce(),
            .sr(N__46911));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_6 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_3_15_6  (
            .in0(N__23036),
            .in1(N__23235),
            .in2(N__19838),
            .in3(N__22617),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47653),
            .ce(),
            .sr(N__46911));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_3_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_3_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_3_15_7 .LUT_INIT=16'b1101110011011000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_3_15_7  (
            .in0(N__22613),
            .in1(N__19829),
            .in2(N__23257),
            .in3(N__23037),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47653),
            .ce(),
            .sr(N__46911));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_3_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_3_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_3_16_0 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_3_16_0  (
            .in0(N__23185),
            .in1(N__23045),
            .in2(N__22608),
            .in3(N__19982),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47642),
            .ce(),
            .sr(N__46916));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_3_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_3_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_3_16_1 .LUT_INIT=16'b1111001111100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_3_16_1  (
            .in0(N__23040),
            .in1(N__22541),
            .in2(N__19976),
            .in3(N__23188),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47642),
            .ce(),
            .sr(N__46916));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_3_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_3_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_3_16_2 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_3_16_2  (
            .in0(N__23183),
            .in1(N__23043),
            .in2(N__22606),
            .in3(N__19967),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47642),
            .ce(),
            .sr(N__46916));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_3_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_3_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_3_16_4 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_3_16_4  (
            .in0(N__23184),
            .in1(N__23044),
            .in2(N__22607),
            .in3(N__19961),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47642),
            .ce(),
            .sr(N__46916));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_3_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_3_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_3_16_5 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_3_16_5  (
            .in0(N__23041),
            .in1(N__23186),
            .in2(N__19955),
            .in3(N__22551),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47642),
            .ce(),
            .sr(N__46916));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_3_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_3_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_3_16_7 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_3_16_7  (
            .in0(N__23042),
            .in1(N__23187),
            .in2(N__19946),
            .in3(N__22552),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47642),
            .ce(),
            .sr(N__46916));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0  (
            .in0(_gnd_net_),
            .in1(N__21638),
            .in2(N__20846),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1  (
            .in0(_gnd_net_),
            .in1(N__22445),
            .in2(N__20885),
            .in3(N__19922),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__47629),
            .ce(),
            .sr(N__46920));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__22454),
            .in2(N__22874),
            .in3(N__19919),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__47629),
            .ce(),
            .sr(N__46920));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__21617),
            .in2(N__22792),
            .in3(N__20051),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__47629),
            .ce(),
            .sr(N__46920));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__22831),
            .in2(N__21677),
            .in3(N__20048),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__47629),
            .ce(),
            .sr(N__46920));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5  (
            .in0(_gnd_net_),
            .in1(N__21263),
            .in2(N__20795),
            .in3(N__20045),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__47629),
            .ce(),
            .sr(N__46920));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__21668),
            .in2(N__22916),
            .in3(N__20042),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__47629),
            .ce(),
            .sr(N__46920));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7  (
            .in0(_gnd_net_),
            .in1(N__21257),
            .in2(N__21251),
            .in3(N__20039),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__47629),
            .ce(),
            .sr(N__46920));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__21650),
            .in2(N__23294),
            .in3(N__20036),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__47618),
            .ce(),
            .sr(N__46925));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__21611),
            .in2(N__21137),
            .in3(N__20024),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__47618),
            .ce(),
            .sr(N__46925));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(N__21656),
            .in2(N__21371),
            .in3(N__20006),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__47618),
            .ce(),
            .sr(N__46925));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3  (
            .in0(_gnd_net_),
            .in1(N__21644),
            .in2(N__21314),
            .in3(N__19985),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__47618),
            .ce(),
            .sr(N__46925));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4  (
            .in0(_gnd_net_),
            .in1(N__21662),
            .in2(N__21167),
            .in3(N__20144),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__47618),
            .ce(),
            .sr(N__46925));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5  (
            .in0(_gnd_net_),
            .in1(N__22008),
            .in2(N__21404),
            .in3(N__20141),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__47618),
            .ce(),
            .sr(N__46925));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6  (
            .in0(_gnd_net_),
            .in1(N__21194),
            .in2(N__22042),
            .in3(N__20123),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__47618),
            .ce(),
            .sr(N__46925));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7  (
            .in0(_gnd_net_),
            .in1(N__22012),
            .in2(N__21101),
            .in3(N__20099),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__47618),
            .ce(),
            .sr(N__46925));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0  (
            .in0(_gnd_net_),
            .in1(N__22013),
            .in2(N__20981),
            .in3(N__20087),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__47606),
            .ce(),
            .sr(N__46929));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__21041),
            .in2(N__22043),
            .in3(N__20075),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__47606),
            .ce(),
            .sr(N__46929));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__22017),
            .in2(N__21068),
            .in3(N__20072),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__47606),
            .ce(),
            .sr(N__46929));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(N__21575),
            .in2(N__22044),
            .in3(N__20069),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__47606),
            .ce(),
            .sr(N__46929));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4  (
            .in0(_gnd_net_),
            .in1(N__22021),
            .in2(N__20954),
            .in3(N__20054),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__47606),
            .ce(),
            .sr(N__46929));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__21011),
            .in2(N__22045),
            .in3(N__20237),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__47606),
            .ce(),
            .sr(N__46929));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6  (
            .in0(_gnd_net_),
            .in1(N__22025),
            .in2(N__22703),
            .in3(N__20222),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__47606),
            .ce(),
            .sr(N__46929));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7  (
            .in0(_gnd_net_),
            .in1(N__21605),
            .in2(N__22046),
            .in3(N__20210),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__47606),
            .ce(),
            .sr(N__46929));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0  (
            .in0(_gnd_net_),
            .in1(N__22029),
            .in2(N__21473),
            .in3(N__20198),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_3_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__47597),
            .ce(),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__21521),
            .in2(N__22047),
            .in3(N__20186),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__47597),
            .ce(),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2  (
            .in0(_gnd_net_),
            .in1(N__22033),
            .in2(N__21440),
            .in3(N__20174),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__47597),
            .ce(),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3  (
            .in0(_gnd_net_),
            .in1(N__21497),
            .in2(N__22048),
            .in3(N__20159),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__47597),
            .ce(),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__22037),
            .in2(N__22742),
            .in3(N__20147),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__47597),
            .ce(),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5  (
            .in0(_gnd_net_),
            .in1(N__21338),
            .in2(N__22049),
            .in3(N__20693),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__47597),
            .ce(),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6  (
            .in0(N__23256),
            .in1(N__22041),
            .in2(_gnd_net_),
            .in3(N__20690),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47597),
            .ce(),
            .sr(N__46932));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_3_21_6  (
            .in0(_gnd_net_),
            .in1(N__20669),
            .in2(_gnd_net_),
            .in3(N__20634),
            .lcout(\current_shift_inst.PI_CTRL.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_21_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_3_21_7  (
            .in0(N__20599),
            .in1(N__20582),
            .in2(N__20567),
            .in3(N__20548),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_22_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_5_LC_3_22_4  (
            .in0(_gnd_net_),
            .in1(N__20520),
            .in2(_gnd_net_),
            .in3(N__20491),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_22_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_3_22_5  (
            .in0(N__20457),
            .in1(N__20425),
            .in2(N__20396),
            .in3(N__20386),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_23_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_23_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_3_23_3  (
            .in0(N__20339),
            .in1(N__20308),
            .in2(N__20285),
            .in3(N__20258),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_3_23_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_3_23_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_3_23_6  (
            .in0(N__23565),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22291),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_3_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_3_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_3_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_3_24_0  (
            .in0(_gnd_net_),
            .in1(N__23530),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_24_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_3_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_3_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_3_24_1  (
            .in0(_gnd_net_),
            .in1(N__20756),
            .in2(_gnd_net_),
            .in3(N__20747),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_3_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_3_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_3_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_3_24_2  (
            .in0(_gnd_net_),
            .in1(N__20744),
            .in2(_gnd_net_),
            .in3(N__20735),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_3_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_3_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_3_24_3  (
            .in0(_gnd_net_),
            .in1(N__20732),
            .in2(_gnd_net_),
            .in3(N__20723),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_3_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_3_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_3_24_4  (
            .in0(_gnd_net_),
            .in1(N__21932),
            .in2(_gnd_net_),
            .in3(N__20720),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_3_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_3_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_3_24_5  (
            .in0(_gnd_net_),
            .in1(N__37818),
            .in2(N__21893),
            .in3(N__20717),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_3_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_3_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_3_24_6  (
            .in0(_gnd_net_),
            .in1(N__21851),
            .in2(N__37917),
            .in3(N__20714),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_3_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_3_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_3_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_3_24_7  (
            .in0(_gnd_net_),
            .in1(N__37822),
            .in2(N__21812),
            .in3(N__20711),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_3_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_3_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_3_25_0  (
            .in0(_gnd_net_),
            .in1(N__21770),
            .in2(_gnd_net_),
            .in3(N__20708),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ),
            .ltout(),
            .carryin(bfn_3_25_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_3_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_3_25_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_3_25_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21731),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_3_25_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_3_25_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_3_25_2  (
            .in0(_gnd_net_),
            .in1(N__21689),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_3_25_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_3_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_3_25_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_3_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22247),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_3_25_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_3_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_3_25_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_3_25_4  (
            .in0(_gnd_net_),
            .in1(N__22202),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_3_25_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_3_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_3_25_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_3_25_5  (
            .in0(_gnd_net_),
            .in1(N__22160),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_3_25_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_3_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_3_25_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_3_25_6  (
            .in0(_gnd_net_),
            .in1(N__22136),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_3_25_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_3_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_3_25_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_3_25_7  (
            .in0(_gnd_net_),
            .in1(N__22112),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_3_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_3_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_3_26_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_3_26_0  (
            .in0(_gnd_net_),
            .in1(N__22088),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_26_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_3_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_3_26_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_3_26_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22064),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_3_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_3_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_3_26_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_3_26_2  (
            .in0(_gnd_net_),
            .in1(N__22337),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_3_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_3_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_3_26_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_3_26_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22325),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_3_26_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_3_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_3_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_3_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20924),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_4_11_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_4_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_4_11_0 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_4_11_0  (
            .in0(N__20921),
            .in1(N__23073),
            .in2(_gnd_net_),
            .in3(N__22612),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47684),
            .ce(),
            .sr(N__46888));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_0 .LUT_INIT=16'b1011000010110001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_4_13_0  (
            .in0(N__22610),
            .in1(N__23261),
            .in2(N__20909),
            .in3(N__23075),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47664),
            .ce(),
            .sr(N__46899));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_4_13_1 .LUT_INIT=16'b1100000011110001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_4_13_1  (
            .in0(N__23074),
            .in1(N__22611),
            .in2(N__20897),
            .in3(N__23260),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47664),
            .ce(),
            .sr(N__46899));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_14_0 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_4_14_0  (
            .in0(N__22873),
            .in1(N__20884),
            .in2(N__20838),
            .in3(N__22791),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_14_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_4_14_1  (
            .in0(N__23283),
            .in1(N__20791),
            .in2(N__20798),
            .in3(N__21218),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_4_14_2  (
            .in0(N__21239),
            .in1(N__20780),
            .in2(N__22908),
            .in3(N__23282),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_14_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_4_14_4  (
            .in0(N__21363),
            .in1(N__21091),
            .in2(N__21313),
            .in3(N__21396),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_14_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_4_14_6  (
            .in0(N__21240),
            .in1(N__22830),
            .in2(_gnd_net_),
            .in3(N__22904),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_4_15_0  (
            .in0(N__21060),
            .in1(N__21036),
            .in2(N__21010),
            .in3(N__20973),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_4_15_1  (
            .in0(N__21186),
            .in1(N__21156),
            .in2(N__21130),
            .in3(N__22732),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_15_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_4_15_2  (
            .in0(N__21212),
            .in1(N__21203),
            .in2(N__21197),
            .in3(N__21533),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_15_3  (
            .in0(N__21185),
            .in1(N__21155),
            .in2(N__21129),
            .in3(N__21089),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_4_15_4  (
            .in0(N__21059),
            .in1(N__21037),
            .in2(N__21009),
            .in3(N__20972),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_4_15_5  (
            .in0(N__23233),
            .in1(N__20946),
            .in2(N__21574),
            .in3(N__21598),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_16_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__21515),
            .in2(_gnd_net_),
            .in3(N__20945),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_16_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_4_16_1  (
            .in0(N__21596),
            .in1(N__21566),
            .in2(N__21545),
            .in3(N__21527),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_16_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_4_16_2  (
            .in0(N__21542),
            .in1(N__23245),
            .in2(N__21536),
            .in3(N__22694),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_16_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_4_16_4  (
            .in0(N__21491),
            .in1(N__21458),
            .in2(N__21439),
            .in3(N__21332),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_4_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_4_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_4_16_5  (
            .in0(N__21516),
            .in1(N__21492),
            .in2(N__21466),
            .in3(N__21435),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__21397),
            .in2(_gnd_net_),
            .in3(N__21364),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_4_16_7  (
            .in0(N__21333),
            .in1(N__21309),
            .in2(N__21272),
            .in3(N__21269),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_4_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_4_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_4_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_4_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25228),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47619),
            .ce(),
            .sr(N__46917));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25159),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47619),
            .ce(),
            .sr(N__46917));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_4_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25261),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47619),
            .ce(),
            .sr(N__46917));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_4_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_4_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25195),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47619),
            .ce(),
            .sr(N__46917));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_4_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25531),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47607),
            .ce(),
            .sr(N__46921));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_4_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_4_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25597),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47607),
            .ce(),
            .sr(N__46921));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_4_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_4_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_4_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25132),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47607),
            .ce(),
            .sr(N__46921));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_4_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_4_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25567),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47607),
            .ce(),
            .sr(N__46921));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_4_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_4_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_4_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_4_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25385),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47607),
            .ce(),
            .sr(N__46921));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_4_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_4_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_4_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_4_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25294),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47607),
            .ce(),
            .sr(N__46921));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_4_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_4_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_4_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_4_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25627),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47598),
            .ce(),
            .sr(N__46926));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_4_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_4_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_4_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_4_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25442),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47598),
            .ce(),
            .sr(N__46926));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_4_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_4_23_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_4_23_0  (
            .in0(_gnd_net_),
            .in1(N__21962),
            .in2(N__21947),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_4_23_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_4_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_4_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_4_23_1  (
            .in0(_gnd_net_),
            .in1(N__21926),
            .in2(N__21908),
            .in3(N__21884),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_4_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_4_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_4_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_4_23_2  (
            .in0(_gnd_net_),
            .in1(N__21881),
            .in2(N__21866),
            .in3(N__21845),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_4_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_4_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_4_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_4_23_3  (
            .in0(_gnd_net_),
            .in1(N__21842),
            .in2(N__21827),
            .in3(N__21803),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_4_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_4_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_4_23_4  (
            .in0(_gnd_net_),
            .in1(N__21800),
            .in2(N__21788),
            .in3(N__21761),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_4_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_4_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_4_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_4_23_5  (
            .in0(_gnd_net_),
            .in1(N__21758),
            .in2(N__21746),
            .in3(N__21719),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_4_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_4_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_4_23_6  (
            .in0(_gnd_net_),
            .in1(N__21716),
            .in2(N__21704),
            .in3(N__21680),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_4_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_4_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_4_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_4_23_7  (
            .in0(_gnd_net_),
            .in1(N__22274),
            .in2(N__22262),
            .in3(N__22235),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_4_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_4_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_4_24_0  (
            .in0(_gnd_net_),
            .in1(N__22232),
            .in2(N__22217),
            .in3(N__22196),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(bfn_4_24_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_4_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_4_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_4_24_1  (
            .in0(_gnd_net_),
            .in1(N__22193),
            .in2(N__22175),
            .in3(N__22154),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_4_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_4_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_4_24_2  (
            .in0(_gnd_net_),
            .in1(N__22151),
            .in2(N__46071),
            .in3(N__22130),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_4_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_4_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_4_24_3  (
            .in0(_gnd_net_),
            .in1(N__22127),
            .in2(N__46073),
            .in3(N__22106),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_4_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_4_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_4_24_4  (
            .in0(_gnd_net_),
            .in1(N__22103),
            .in2(N__46072),
            .in3(N__22079),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_4_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_4_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_4_24_5  (
            .in0(_gnd_net_),
            .in1(N__22076),
            .in2(N__46074),
            .in3(N__22052),
            .lcout(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_4_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_4_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_4_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_4_24_6  (
            .in0(_gnd_net_),
            .in1(N__46064),
            .in2(N__22352),
            .in3(N__22328),
            .lcout(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_4_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_4_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_4_24_7  (
            .in0(_gnd_net_),
            .in1(N__46057),
            .in2(N__46010),
            .in3(N__22313),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_4_25_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_4_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_4_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_4_25_0  (
            .in0(N__23456),
            .in1(N__22310),
            .in2(_gnd_net_),
            .in3(N__22304),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ),
            .ltout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_1 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_1  (
            .in0(N__23801),
            .in1(N__22420),
            .in2(N__22301),
            .in3(N__23818),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_4_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_4_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_4_25_2 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_4_25_2  (
            .in0(N__23741),
            .in1(N__23758),
            .in2(N__22385),
            .in3(N__24011),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_4 .LUT_INIT=16'b1100001110101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_4  (
            .in0(N__23419),
            .in1(N__23768),
            .in2(N__23792),
            .in3(N__24010),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_4_25_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_4_25_5 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_4_25_5  (
            .in0(N__23693),
            .in1(N__22399),
            .in2(N__24030),
            .in3(N__23710),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_6  (
            .in0(N__23543),
            .in1(N__23569),
            .in2(N__22298),
            .in3(N__24009),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_4_26_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_4_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_4_26_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_4_26_0  (
            .in0(_gnd_net_),
            .in1(N__22435),
            .in2(_gnd_net_),
            .in3(N__23732),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(\pwm_generator_inst.un15_threshold_1_axb_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_4_26_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_4_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_4_26_1 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_4_26_1  (
            .in0(N__22436),
            .in1(N__24019),
            .in2(N__22424),
            .in3(N__23720),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_4_26_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_4_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_4_26_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_4_26_2  (
            .in0(N__23509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23443),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_26_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_26_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_26_3  (
            .in0(_gnd_net_),
            .in1(N__22421),
            .in2(_gnd_net_),
            .in3(N__23819),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_4_26_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_4_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_4_26_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_4_26_5  (
            .in0(N__22400),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23711),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_4_26_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_4_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_4_26_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_4_26_6  (
            .in0(_gnd_net_),
            .in1(N__22384),
            .in2(_gnd_net_),
            .in3(N__23759),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_4_26_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_4_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_4_26_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_4_26_7  (
            .in0(_gnd_net_),
            .in1(N__24079),
            .in2(_gnd_net_),
            .in3(N__24100),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_LC_5_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_5_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_5_10_7 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_5_10_7  (
            .in0(N__23918),
            .in1(N__24913),
            .in2(N__22367),
            .in3(N__32368),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47685),
            .ce(),
            .sr(N__46878));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_5_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_5_11_3 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_5_11_3  (
            .in0(N__23915),
            .in1(N__22363),
            .in2(_gnd_net_),
            .in3(N__33763),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_5_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_5_11_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_5_11_7  (
            .in0(N__23916),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33764),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_5_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_5_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_5_12_4 .LUT_INIT=16'b1011101000001010;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_5_12_4  (
            .in0(N__34588),
            .in1(N__24914),
            .in2(N__32377),
            .in3(N__23917),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47665),
            .ce(),
            .sr(N__46889));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_5_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_5_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_5_14_1 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_5_14_1  (
            .in0(N__23253),
            .in1(N__23050),
            .in2(N__23306),
            .in3(N__22565),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47643),
            .ce(),
            .sr(N__46900));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_7 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_5_14_7  (
            .in0(N__23252),
            .in1(N__23049),
            .in2(N__22931),
            .in3(N__22564),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47643),
            .ce(),
            .sr(N__46900));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_15_5 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_5_15_5  (
            .in0(N__22869),
            .in1(N__22832),
            .in2(N__22793),
            .in3(N__22748),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_5_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_5_15_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_5_15_6  (
            .in0(N__22731),
            .in1(N__22699),
            .in2(N__22670),
            .in3(N__22667),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_16_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_16_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_16_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_5_16_7  (
            .in0(N__22661),
            .in1(N__22655),
            .in2(N__22649),
            .in3(N__22640),
            .lcout(\current_shift_inst.PI_CTRL.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_5_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25324),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47608),
            .ce(),
            .sr(N__46912));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_5_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25354),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47608),
            .ce(),
            .sr(N__46912));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_5_23_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_5_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_5_23_4 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_5_23_4  (
            .in0(N__46283),
            .in1(N__23477),
            .in2(N__46208),
            .in3(N__46075),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_5_24_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_5_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_5_24_5 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_5_24_5  (
            .in0(N__23489),
            .in1(N__23510),
            .in2(N__23444),
            .in3(N__24018),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_5_24_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_5_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_5_24_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_5_24_7  (
            .in0(_gnd_net_),
            .in1(N__23420),
            .in2(_gnd_net_),
            .in3(N__23790),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_5_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_5_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_5_25_0  (
            .in0(_gnd_net_),
            .in1(N__23390),
            .in2(_gnd_net_),
            .in3(N__23405),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_5_25_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_5_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_5_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_5_25_1  (
            .in0(_gnd_net_),
            .in1(N__23369),
            .in2(_gnd_net_),
            .in3(N__23384),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_5_25_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_5_25_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_5_25_2  (
            .in0(_gnd_net_),
            .in1(N__23351),
            .in2(_gnd_net_),
            .in3(N__23363),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_5_25_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_5_25_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_5_25_3  (
            .in0(_gnd_net_),
            .in1(N__23333),
            .in2(_gnd_net_),
            .in3(N__23345),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_5_25_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_5_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_5_25_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_5_25_4  (
            .in0(_gnd_net_),
            .in1(N__23312),
            .in2(_gnd_net_),
            .in3(N__23327),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_5_25_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_5_25_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_5_25_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_5_25_5  (
            .in0(_gnd_net_),
            .in1(N__23660),
            .in2(_gnd_net_),
            .in3(N__23675),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_5_25_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_5_25_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_5_25_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_5_25_6  (
            .in0(_gnd_net_),
            .in1(N__23639),
            .in2(_gnd_net_),
            .in3(N__23654),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_5_25_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_5_25_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_5_25_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_5_25_7  (
            .in0(_gnd_net_),
            .in1(N__23618),
            .in2(_gnd_net_),
            .in3(N__23633),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_5_26_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_5_26_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_5_26_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_5_26_0  (
            .in0(_gnd_net_),
            .in1(N__23597),
            .in2(_gnd_net_),
            .in3(N__23612),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_5_26_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_5_26_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_5_26_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_5_26_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_5_26_1  (
            .in0(_gnd_net_),
            .in1(N__23576),
            .in2(_gnd_net_),
            .in3(N__23591),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_5_26_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_5_26_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_5_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_5_26_2  (
            .in0(_gnd_net_),
            .in1(N__23570),
            .in2(_gnd_net_),
            .in3(N__23537),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_5_26_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_5_26_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_5_26_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_5_26_3  (
            .in0(N__24031),
            .in1(N__23534),
            .in2(_gnd_net_),
            .in3(N__23513),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_5_26_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_5_26_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_5_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_5_26_4  (
            .in0(_gnd_net_),
            .in1(N__23505),
            .in2(_gnd_net_),
            .in3(N__23480),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_5_26_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_5_26_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_5_26_5  (
            .in0(_gnd_net_),
            .in1(N__23817),
            .in2(_gnd_net_),
            .in3(N__23795),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_5_26_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_5_26_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_5_26_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_5_26_6  (
            .in0(_gnd_net_),
            .in1(N__23791),
            .in2(_gnd_net_),
            .in3(N__23762),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_5_26_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_5_26_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_5_26_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_5_26_7  (
            .in0(_gnd_net_),
            .in1(N__23757),
            .in2(_gnd_net_),
            .in3(N__23735),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_5_27_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_5_27_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_5_27_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_5_27_0  (
            .in0(_gnd_net_),
            .in1(N__23731),
            .in2(_gnd_net_),
            .in3(N__23714),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_5_27_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_5_27_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_5_27_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_5_27_1  (
            .in0(_gnd_net_),
            .in1(N__23709),
            .in2(_gnd_net_),
            .in3(N__23684),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_5_27_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_5_27_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_5_27_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_5_27_2  (
            .in0(_gnd_net_),
            .in1(N__24099),
            .in2(_gnd_net_),
            .in3(N__23681),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_5_27_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_5_27_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_5_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_5_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23678),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_7_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_7_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_7_6_4  (
            .in0(N__27207),
            .in1(N__29008),
            .in2(_gnd_net_),
            .in3(N__31993),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_7_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_7_7_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_7_7_4  (
            .in0(N__26980),
            .in1(N__31989),
            .in2(_gnd_net_),
            .in3(N__26960),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_7_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_7_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_7_7_5  (
            .in0(N__31992),
            .in1(N__26100),
            .in2(_gnd_net_),
            .in3(N__26077),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_7_7_6  (
            .in0(N__26041),
            .in1(N__27751),
            .in2(_gnd_net_),
            .in3(N__31991),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_7_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_7_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_7_7_7  (
            .in0(N__31990),
            .in1(N__26184),
            .in2(_gnd_net_),
            .in3(N__27683),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_7_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_7_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_7_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_25_LC_7_8_1  (
            .in0(N__27208),
            .in1(N__29007),
            .in2(_gnd_net_),
            .in3(N__31995),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47686),
            .ce(N__32574),
            .sr(N__46859));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_7_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_7_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_7_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_7_8_3  (
            .in0(N__26958),
            .in1(N__26976),
            .in2(_gnd_net_),
            .in3(N__31994),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47686),
            .ce(N__32574),
            .sr(N__46859));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_7_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_7_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_7_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_7_8_7  (
            .in0(N__26037),
            .in1(N__27752),
            .in2(_gnd_net_),
            .in3(N__31996),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47686),
            .ce(N__32574),
            .sr(N__46859));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_7_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_7_9_1 .LUT_INIT=16'b1111011100110001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_7_9_1  (
            .in0(N__24346),
            .in1(N__24315),
            .in2(N__25019),
            .in3(N__23953),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_7_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_7_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_7_9_3  (
            .in0(N__27607),
            .in1(N__31939),
            .in2(_gnd_net_),
            .in3(N__26014),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(elapsed_time_ns_1_RNIH33T9_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_7_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_7_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_7_9_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_7_9_4  (
            .in0(N__31940),
            .in1(_gnd_net_),
            .in2(N__23822),
            .in3(N__27608),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47675),
            .ce(N__32654),
            .sr(N__46864));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_7_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_7_10_0 .LUT_INIT=16'b0111001100010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_7_10_0  (
            .in0(N__24403),
            .in1(N__24379),
            .in2(N__25034),
            .in3(N__23837),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_7_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_7_10_1 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_7_10_1  (
            .in0(N__23836),
            .in1(N__24404),
            .in2(N__24383),
            .in3(N__25030),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_7_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_7_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_21_LC_7_10_3  (
            .in0(N__31941),
            .in1(N__31453),
            .in2(_gnd_net_),
            .in3(N__31420),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47666),
            .ce(N__32655),
            .sr(N__46869));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_7_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_7_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_7_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_7_10_7  (
            .in0(N__31942),
            .in1(N__26102),
            .in2(_gnd_net_),
            .in3(N__26073),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47666),
            .ce(N__32655),
            .sr(N__46869));
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_7_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_7_11_1 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_RNIO0241_0_30_LC_7_11_1  (
            .in0(N__26331),
            .in1(N__24513),
            .in2(N__23940),
            .in3(N__24540),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_7_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_7_11_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3_28_LC_7_11_2  (
            .in0(N__32373),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32395),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIP2UJ3Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_7_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_7_11_3 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_RNIO0241_30_LC_7_11_3  (
            .in0(N__26332),
            .in1(N__24514),
            .in2(N__23941),
            .in3(N__24541),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un4_running_df30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_7_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_7_11_4 .LUT_INIT=16'b1111110101011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI4E6P2_28_LC_7_11_4  (
            .in0(N__23903),
            .in1(N__24937),
            .in2(N__23828),
            .in3(N__24926),
            .lcout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23825),
            .in3(N__32372),
            .lcout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_7_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_7_11_7 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_7_11_7  (
            .in0(N__26333),
            .in1(N__24515),
            .in2(N__23942),
            .in3(N__24542),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_7_12_0  (
            .in0(N__26945),
            .in1(N__27735),
            .in2(N__27677),
            .in3(N__26060),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_7_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_7_12_5 .LUT_INIT=16'b0100111100000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_7_12_5  (
            .in0(N__24350),
            .in1(N__25012),
            .in2(N__24323),
            .in3(N__23957),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_7_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_7_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_31_LC_7_13_4  (
            .in0(N__28718),
            .in1(N__27817),
            .in2(_gnd_net_),
            .in3(N__31959),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47630),
            .ce(N__32653),
            .sr(N__46884));
    defparam \phase_controller_inst1.state_4_LC_7_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_7_15_2 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_7_15_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.state_4_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__30811),
            .in2(_gnd_net_),
            .in3(N__34661),
            .lcout(phase_controller_inst1_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47609),
            .ce(),
            .sr(N__46894));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_7_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_7_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_7_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33762),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47590),
            .ce(),
            .sr(N__46904));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_17_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_7_17_7 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_7_17_7  (
            .in0(N__29277),
            .in1(N__32963),
            .in2(_gnd_net_),
            .in3(N__30920),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47590),
            .ce(),
            .sr(N__46904));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_7_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_7_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__23879),
            .in2(N__24054),
            .in3(N__24053),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ),
            .ltout(),
            .carryin(bfn_7_23_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_7_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_7_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_7_23_1  (
            .in0(_gnd_net_),
            .in1(N__23867),
            .in2(_gnd_net_),
            .in3(N__23855),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_7_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_7_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_7_23_2  (
            .in0(_gnd_net_),
            .in1(N__23852),
            .in2(_gnd_net_),
            .in3(N__23840),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_7_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_7_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_7_23_3  (
            .in0(_gnd_net_),
            .in1(N__24209),
            .in2(_gnd_net_),
            .in3(N__24197),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_7_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_7_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_7_23_4  (
            .in0(_gnd_net_),
            .in1(N__24194),
            .in2(_gnd_net_),
            .in3(N__24182),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_7_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_7_23_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_7_23_5  (
            .in0(_gnd_net_),
            .in1(N__24179),
            .in2(_gnd_net_),
            .in3(N__24167),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_7_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_7_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_7_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_7_23_6  (
            .in0(_gnd_net_),
            .in1(N__24164),
            .in2(_gnd_net_),
            .in3(N__24152),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_7_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_7_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_7_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_7_23_7  (
            .in0(_gnd_net_),
            .in1(N__24149),
            .in2(_gnd_net_),
            .in3(N__24137),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_7_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_7_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_7_24_0  (
            .in0(_gnd_net_),
            .in1(N__23963),
            .in2(_gnd_net_),
            .in3(N__24134),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ),
            .ltout(),
            .carryin(bfn_7_24_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_7_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_7_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_7_24_1 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_7_24_1  (
            .in0(N__24131),
            .in1(N__24119),
            .in2(N__24056),
            .in3(N__24107),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_7_25_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_7_25_3 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_7_25_3  (
            .in0(N__24104),
            .in1(N__24080),
            .in2(N__24055),
            .in3(N__23975),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D1_LC_8_3_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MAX_D1_LC_8_3_1 (
            .in0(N__24266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_max_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47702),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_4_4 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_8_4_4  (
            .in0(N__25954),
            .in1(N__25903),
            .in2(N__25931),
            .in3(N__25888),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__24257),
            .in2(N__32342),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_8_5_1  (
            .in0(N__32659),
            .in1(N__24469),
            .in2(_gnd_net_),
            .in3(N__24242),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__47698),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_5_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_8_5_2  (
            .in0(N__32598),
            .in1(N__24439),
            .in2(N__24239),
            .in3(N__24224),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__47698),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_8_5_3  (
            .in0(N__32660),
            .in1(N__24724),
            .in2(_gnd_net_),
            .in3(N__24221),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__47698),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_8_5_4  (
            .in0(N__32599),
            .in1(N__24700),
            .in2(_gnd_net_),
            .in3(N__24218),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__47698),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_8_5_5  (
            .in0(N__32661),
            .in1(N__24670),
            .in2(_gnd_net_),
            .in3(N__24215),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__47698),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_8_5_6  (
            .in0(N__32600),
            .in1(N__24649),
            .in2(_gnd_net_),
            .in3(N__24212),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__47698),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_8_5_7  (
            .in0(N__32662),
            .in1(N__24625),
            .in2(_gnd_net_),
            .in3(N__24293),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__47698),
            .ce(),
            .sr(N__46835));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_8_6_0  (
            .in0(N__32670),
            .in1(N__24601),
            .in2(_gnd_net_),
            .in3(N__24290),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__47695),
            .ce(),
            .sr(N__46842));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_8_6_1  (
            .in0(N__32609),
            .in1(N__24577),
            .in2(_gnd_net_),
            .in3(N__24287),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__47695),
            .ce(),
            .sr(N__46842));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_8_6_2  (
            .in0(N__32667),
            .in1(N__24880),
            .in2(_gnd_net_),
            .in3(N__24284),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__47695),
            .ce(),
            .sr(N__46842));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_8_6_3  (
            .in0(N__32610),
            .in1(N__24853),
            .in2(_gnd_net_),
            .in3(N__24281),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__47695),
            .ce(),
            .sr(N__46842));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_8_6_4  (
            .in0(N__32668),
            .in1(N__24829),
            .in2(_gnd_net_),
            .in3(N__24278),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__47695),
            .ce(),
            .sr(N__46842));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_8_6_5  (
            .in0(N__32611),
            .in1(N__24802),
            .in2(_gnd_net_),
            .in3(N__24275),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__47695),
            .ce(),
            .sr(N__46842));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_8_6_6  (
            .in0(N__32669),
            .in1(N__24781),
            .in2(_gnd_net_),
            .in3(N__24272),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__47695),
            .ce(),
            .sr(N__46842));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_8_6_7  (
            .in0(N__32612),
            .in1(N__25927),
            .in2(_gnd_net_),
            .in3(N__24269),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__47695),
            .ce(),
            .sr(N__46842));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_8_7_0  (
            .in0(N__32605),
            .in1(N__25953),
            .in2(_gnd_net_),
            .in3(N__24413),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__47687),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_8_7_1  (
            .in0(N__32663),
            .in1(N__25823),
            .in2(_gnd_net_),
            .in3(N__24410),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__47687),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_8_7_2  (
            .in0(N__32606),
            .in1(N__25838),
            .in2(_gnd_net_),
            .in3(N__24407),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__47687),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_8_7_3  (
            .in0(N__32664),
            .in1(N__24402),
            .in2(_gnd_net_),
            .in3(N__24386),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__47687),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_8_7_4  (
            .in0(N__32607),
            .in1(N__24373),
            .in2(_gnd_net_),
            .in3(N__24359),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__47687),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_8_7_5  (
            .in0(N__32665),
            .in1(N__25970),
            .in2(_gnd_net_),
            .in3(N__24356),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__47687),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_8_7_6  (
            .in0(N__32608),
            .in1(N__25987),
            .in2(_gnd_net_),
            .in3(N__24353),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__47687),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_8_7_7  (
            .in0(N__32666),
            .in1(N__24345),
            .in2(_gnd_net_),
            .in3(N__24326),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__47687),
            .ce(),
            .sr(N__46847));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_8_8_0  (
            .in0(N__32552),
            .in1(N__24316),
            .in2(_gnd_net_),
            .in3(N__24296),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__47676),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_8_8_1  (
            .in0(N__32571),
            .in1(N__25071),
            .in2(_gnd_net_),
            .in3(N__24554),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__47676),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_8_8_2  (
            .in0(N__32553),
            .in1(N__25092),
            .in2(_gnd_net_),
            .in3(N__24551),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__47676),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_8_8_3  (
            .in0(N__32572),
            .in1(N__30981),
            .in2(_gnd_net_),
            .in3(N__24548),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__47676),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_8_8_4  (
            .in0(N__32554),
            .in1(N__30957),
            .in2(_gnd_net_),
            .in3(N__24545),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__47676),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_8_8_5  (
            .in0(N__32573),
            .in1(N__24539),
            .in2(_gnd_net_),
            .in3(N__24521),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__47676),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_8_8_6  (
            .in0(N__32555),
            .in1(N__24512),
            .in2(_gnd_net_),
            .in3(N__24518),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47676),
            .ce(),
            .sr(N__46853));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_8_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_8_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__24491),
            .in2(N__24485),
            .in3(N__32335),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_8_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_8_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__24476),
            .in2(N__24455),
            .in3(N__24470),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_8_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_8_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__24446),
            .in2(N__24425),
            .in3(N__24440),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_8_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_8_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__26165),
            .in2(N__24710),
            .in3(N__24728),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_8_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_8_9_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_8_9_4  (
            .in0(N__24701),
            .in1(N__24677),
            .in2(N__24686),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_8_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_8_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_8_9_5  (
            .in0(N__24671),
            .in1(N__24656),
            .in2(N__26300),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_8_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_8_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_8_9_6  (
            .in0(N__24650),
            .in1(N__31532),
            .in2(N__24635),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_8_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_8_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_8_9_7  (
            .in0(N__24626),
            .in1(N__25046),
            .in2(N__24611),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_8_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_8_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_8_10_0  (
            .in0(N__24602),
            .in1(N__26234),
            .in2(N__24587),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_8_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_8_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__26249),
            .in2(N__24563),
            .in3(N__24578),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_8_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_8_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__26339),
            .in2(N__24866),
            .in3(N__24881),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_8_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_8_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__26285),
            .in2(N__24839),
            .in3(N__24857),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_8_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_8_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__26315),
            .in2(N__24815),
            .in3(N__24830),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_8_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_8_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_8_10_5  (
            .in0(N__24803),
            .in1(N__24788),
            .in2(N__27041),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_8_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_8_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_8_10_6  (
            .in0(N__24782),
            .in1(N__25790),
            .in2(N__24767),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_8_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_8_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__24755),
            .in2(N__25877),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_8_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__25862),
            .in2(N__25808),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_8_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_8_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__24743),
            .in2(N__24737),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_8_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_8_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__26228),
            .in2(N__26003),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_8_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_8_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__24968),
            .in2(N__24962),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_8_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_8_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__24887),
            .in2(N__25055),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_8_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_8_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__30932),
            .in2(N__31064),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_8_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_8_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__24950),
            .in2(N__24944),
            .in3(N__24920),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_8_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_8_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24917),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_8_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_8_12_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_8_12_2  (
            .in0(N__28903),
            .in1(N__31764),
            .in2(_gnd_net_),
            .in3(N__27391),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(elapsed_time_ns_1_RNI58DN9_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_8_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_8_12_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_27_LC_8_12_3  (
            .in0(N__31765),
            .in1(_gnd_net_),
            .in2(N__24890),
            .in3(N__28904),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47631),
            .ce(N__32647),
            .sr(N__46873));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_8_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_8_12_4 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_8_12_4  (
            .in0(N__26308),
            .in1(N__25093),
            .in2(N__25076),
            .in3(N__25105),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_8_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_8_12_5 .LUT_INIT=16'b0000101010001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_8_12_5  (
            .in0(N__25106),
            .in1(N__26309),
            .in2(N__25097),
            .in3(N__25075),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_8_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_8_13_1  (
            .in0(N__31770),
            .in1(N__29424),
            .in2(_gnd_net_),
            .in3(N__29408),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47620),
            .ce(N__32652),
            .sr(N__46879));
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_8_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_8_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_8_13_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_20_LC_8_13_2  (
            .in0(N__31565),
            .in1(N__32040),
            .in2(_gnd_net_),
            .in3(N__31771),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47620),
            .ce(N__32652),
            .sr(N__46879));
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_8_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_8_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_24_LC_8_13_5  (
            .in0(N__31769),
            .in1(N__26913),
            .in2(_gnd_net_),
            .in3(N__29075),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47620),
            .ce(N__32652),
            .sr(N__46879));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_14_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27772),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47610),
            .ce(N__28683),
            .sr(N__46885));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_15_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27703),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47599),
            .ce(N__28671),
            .sr(N__46890));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_16_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(N__29276),
            .in2(_gnd_net_),
            .in3(N__30919),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_202_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__29126),
            .in2(_gnd_net_),
            .in3(N__29300),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47584),
            .ce(),
            .sr(N__46901));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_8_19_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_8_19_0  (
            .in0(N__26504),
            .in1(N__24974),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_8_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_8_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__26498),
            .in2(_gnd_net_),
            .in3(N__25358),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__47574),
            .ce(),
            .sr(N__46908));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_8_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_8_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__26489),
            .in2(_gnd_net_),
            .in3(N__25328),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__47574),
            .ce(),
            .sr(N__46908));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_8_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_8_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__26594),
            .in2(_gnd_net_),
            .in3(N__25298),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__47574),
            .ce(),
            .sr(N__46908));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_8_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_8_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__26585),
            .in2(_gnd_net_),
            .in3(N__25268),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__47574),
            .ce(),
            .sr(N__46908));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_8_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_8_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__26576),
            .in2(_gnd_net_),
            .in3(N__25235),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__47574),
            .ce(),
            .sr(N__46908));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_8_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__26567),
            .in2(_gnd_net_),
            .in3(N__25202),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__47574),
            .ce(),
            .sr(N__46908));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_8_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_8_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__26558),
            .in2(_gnd_net_),
            .in3(N__25169),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__47574),
            .ce(),
            .sr(N__46908));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_8_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_8_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__26549),
            .in2(_gnd_net_),
            .in3(N__25139),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__47569),
            .ce(),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_8_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_8_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_8_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__26540),
            .in2(_gnd_net_),
            .in3(N__25634),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__47569),
            .ce(),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_8_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_8_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_8_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__26531),
            .in2(_gnd_net_),
            .in3(N__25601),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__47569),
            .ce(),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_8_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_8_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__26708),
            .in2(_gnd_net_),
            .in3(N__25571),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__47569),
            .ce(),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_8_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_8_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_8_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__26699),
            .in2(_gnd_net_),
            .in3(N__25541),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__47569),
            .ce(),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_8_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_8_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_8_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_8_20_5  (
            .in0(_gnd_net_),
            .in1(N__26675),
            .in2(_gnd_net_),
            .in3(N__25505),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__47569),
            .ce(),
            .sr(N__46913));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_8_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_8_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_8_20_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(N__26687),
            .in2(_gnd_net_),
            .in3(N__25502),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47569),
            .ce(),
            .sr(N__46913));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_8_23_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_8_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_8_23_1 .LUT_INIT=16'b1111001111110101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_8_23_1  (
            .in0(N__25690),
            .in1(N__25735),
            .in2(N__25412),
            .in3(N__46169),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_8_23_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_8_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_8_23_2 .LUT_INIT=16'b1111010111110011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_8_23_2  (
            .in0(N__25736),
            .in1(N__25691),
            .in2(N__25403),
            .in3(N__46249),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_8_23_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_8_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_8_23_4 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_8_23_4  (
            .in0(N__25734),
            .in1(N__25689),
            .in2(N__25394),
            .in3(N__46248),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_8_23_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_8_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_8_23_6 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_8_23_6  (
            .in0(N__25733),
            .in1(N__25688),
            .in2(N__25778),
            .in3(N__46247),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_8_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_8_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_8_23_7 .LUT_INIT=16'b1100110111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_8_23_7  (
            .in0(N__25687),
            .in1(N__25769),
            .in2(N__46255),
            .in3(N__25732),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_8_24_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_8_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_8_24_0 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_8_24_0  (
            .in0(N__25719),
            .in1(N__25685),
            .in2(N__46259),
            .in3(N__25763),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_8_24_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_8_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_8_24_2 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_8_24_2  (
            .in0(N__25720),
            .in1(N__46243),
            .in2(N__25757),
            .in3(N__25686),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_8_24_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_8_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_8_24_3 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_8_24_3  (
            .in0(N__25684),
            .in1(N__25748),
            .in2(N__46254),
            .in3(N__25718),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_24_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_24_5 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_24_5  (
            .in0(N__25682),
            .in1(N__25742),
            .in2(N__46253),
            .in3(N__25716),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_8_24_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_8_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_8_24_6 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_8_24_6  (
            .in0(N__25717),
            .in1(N__25683),
            .in2(N__25643),
            .in3(N__46242),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_3_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_3_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_9_3_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_9_3_5  (
            .in0(N__29730),
            .in1(N__29713),
            .in2(_gnd_net_),
            .in3(N__31911),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47701),
            .ce(N__32657),
            .sr(N__46812));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_4_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_9_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_9_4_0  (
            .in0(N__26895),
            .in1(N__28571),
            .in2(_gnd_net_),
            .in3(N__32009),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47699),
            .ce(N__32658),
            .sr(N__46821));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_5_0 .LUT_INIT=16'b0111010100010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_9_5_0  (
            .in0(N__25955),
            .in1(N__25926),
            .in2(N__25907),
            .in3(N__25889),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_9_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_9_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_9_5_2  (
            .in0(N__31969),
            .in1(N__26897),
            .in2(_gnd_net_),
            .in3(N__28569),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_9_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_9_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_9_5_5  (
            .in0(N__26851),
            .in1(N__27910),
            .in2(_gnd_net_),
            .in3(N__31968),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_6_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_6_0  (
            .in0(N__25847),
            .in1(N__25837),
            .in2(N__27059),
            .in3(N__25822),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_9_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_9_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_9_6_1  (
            .in0(N__31965),
            .in1(N__28503),
            .in2(_gnd_net_),
            .in3(N__27004),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(elapsed_time_ns_1_RNI57CN9_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_9_6_2 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_9_6_2  (
            .in0(N__28504),
            .in1(N__31967),
            .in2(N__25850),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47688),
            .ce(N__32671),
            .sr(N__46836));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_6_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_9_6_4  (
            .in0(N__25846),
            .in1(N__25836),
            .in2(N__27058),
            .in3(N__25821),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_6_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_9_6_5  (
            .in0(N__31963),
            .in1(N__29619),
            .in2(_gnd_net_),
            .in3(N__29584),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(elapsed_time_ns_1_RNI24CN9_0_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_9_6_6 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_9_6_6  (
            .in0(N__29620),
            .in1(N__31966),
            .in2(N__25793),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47688),
            .ce(N__32671),
            .sr(N__46836));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_9_6_7  (
            .in0(N__31964),
            .in1(N__27079),
            .in2(_gnd_net_),
            .in3(N__28435),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_9_7_0  (
            .in0(N__30115),
            .in1(N__26993),
            .in2(N__26114),
            .in3(N__30415),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_9_7_1  (
            .in0(N__26992),
            .in1(N__30116),
            .in2(N__30419),
            .in3(N__26110),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_9_7_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_9_7_3  (
            .in0(N__27075),
            .in1(N__31972),
            .in2(_gnd_net_),
            .in3(N__28433),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__31312),
            .sr(N__46843));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_9_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_9_7_4  (
            .in0(N__31970),
            .in1(N__26101),
            .in2(_gnd_net_),
            .in3(N__26078),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__31312),
            .sr(N__46843));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_9_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_9_7_5  (
            .in0(N__26042),
            .in1(N__31973),
            .in2(_gnd_net_),
            .in3(N__27750),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__31312),
            .sr(N__46843));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_9_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_9_7_6  (
            .in0(N__31971),
            .in1(N__26185),
            .in2(_gnd_net_),
            .in3(N__27681),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__31312),
            .sr(N__46843));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_9_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_9_7_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_9_7_7  (
            .in0(N__27606),
            .in1(N__31974),
            .in2(_gnd_net_),
            .in3(N__26021),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47677),
            .ce(N__31312),
            .sr(N__46843));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_8_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_8_0  (
            .in0(N__25969),
            .in1(N__26198),
            .in2(N__26213),
            .in3(N__25986),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_8_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_9_8_1  (
            .in0(N__26197),
            .in1(N__26209),
            .in2(N__25988),
            .in3(N__25968),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_9_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_9_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_9_8_2  (
            .in0(N__28248),
            .in1(N__26137),
            .in2(_gnd_net_),
            .in3(N__31907),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(elapsed_time_ns_1_RNI14DN9_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_9_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_9_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_9_8_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_23_LC_9_8_3  (
            .in0(N__31909),
            .in1(_gnd_net_),
            .in2(N__26216),
            .in3(N__28249),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47667),
            .ce(N__32601),
            .sr(N__46848));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_9_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_9_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_9_8_4  (
            .in0(N__28305),
            .in1(N__31906),
            .in2(_gnd_net_),
            .in3(N__26158),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(elapsed_time_ns_1_RNI03DN9_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_9_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_9_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_9_8_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_22_LC_9_8_5  (
            .in0(N__31908),
            .in1(_gnd_net_),
            .in2(N__26201),
            .in3(N__28306),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47667),
            .ce(N__32601),
            .sr(N__46848));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_9_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_9_8_7  (
            .in0(N__31910),
            .in1(N__26189),
            .in2(_gnd_net_),
            .in3(N__27682),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47667),
            .ce(N__32601),
            .sr(N__46848));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_9_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_9_9_0  (
            .in0(N__30359),
            .in1(N__30382),
            .in2(N__26126),
            .in3(N__26147),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_9_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_9_9_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_9_9_1  (
            .in0(N__26146),
            .in1(N__30358),
            .in2(N__30386),
            .in3(N__26122),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_9_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_9_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_22_LC_9_9_2  (
            .in0(N__31901),
            .in1(N__28307),
            .in2(_gnd_net_),
            .in3(N__26159),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47654),
            .ce(N__31311),
            .sr(N__46854));
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_9_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_9_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_23_LC_9_9_3  (
            .in0(N__26138),
            .in1(N__28250),
            .in2(_gnd_net_),
            .in3(N__31903),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47654),
            .ce(N__31311),
            .sr(N__46854));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_9_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_9_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_9_9_6  (
            .in0(N__31900),
            .in1(N__26363),
            .in2(_gnd_net_),
            .in3(N__28049),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47654),
            .ce(N__31311),
            .sr(N__46854));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_9_9_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_9_9_7  (
            .in0(N__28112),
            .in1(N__31902),
            .in2(_gnd_net_),
            .in3(N__26264),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47654),
            .ce(N__31311),
            .sr(N__46854));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_9_10_0  (
            .in0(N__28154),
            .in1(N__27981),
            .in2(N__28111),
            .in3(N__28044),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_9_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_9_10_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_9_10_1  (
            .in0(N__27597),
            .in1(N__27550),
            .in2(N__26267),
            .in3(N__26243),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_9_10_2  (
            .in0(N__28106),
            .in1(_gnd_net_),
            .in2(N__31988),
            .in3(N__26263),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(elapsed_time_ns_1_RNITUBN9_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_9_10_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__28107),
            .in2(N__26252),
            .in3(N__31898),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__32616),
            .sr(N__46860));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_9_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_9_10_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__29400),
            .in2(_gnd_net_),
            .in3(N__31362),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_9_10_5  (
            .in0(N__27019),
            .in1(N__31894),
            .in2(_gnd_net_),
            .in3(N__28155),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(elapsed_time_ns_1_RNIL73T9_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_9_10_6  (
            .in0(N__28156),
            .in1(_gnd_net_),
            .in2(N__26237),
            .in3(N__31912),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__32616),
            .sr(N__46860));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_9_10_7  (
            .in0(N__28045),
            .in1(N__26359),
            .in2(_gnd_net_),
            .in3(N__31899),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47644),
            .ce(N__32616),
            .sr(N__46860));
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_9_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_9_11_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_30_LC_9_11_0  (
            .in0(N__27789),
            .in1(N__28760),
            .in2(_gnd_net_),
            .in3(N__31779),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47632),
            .ce(N__32590),
            .sr(N__46865));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_9_11_1  (
            .in0(N__30470),
            .in1(N__31904),
            .in2(_gnd_net_),
            .in3(N__30443),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47632),
            .ce(N__32590),
            .sr(N__46865));
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_9_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_9_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_9_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_26_LC_9_11_2  (
            .in0(N__30749),
            .in1(N__30779),
            .in2(_gnd_net_),
            .in3(N__31778),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47632),
            .ce(N__32590),
            .sr(N__46865));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_9_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_9_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_9_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_9_11_4  (
            .in0(N__27549),
            .in1(N__26871),
            .in2(_gnd_net_),
            .in3(N__31780),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47632),
            .ce(N__32590),
            .sr(N__46865));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_9_11_6  (
            .in0(N__27441),
            .in1(N__27983),
            .in2(_gnd_net_),
            .in3(N__31777),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47632),
            .ce(N__32590),
            .sr(N__46865));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_9_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_9_12_0 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_9_12_0  (
            .in0(N__28709),
            .in1(N__26279),
            .in2(N__26372),
            .in3(N__26387),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_9_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_9_12_1 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_9_12_1  (
            .in0(N__31446),
            .in1(_gnd_net_),
            .in2(N__26270),
            .in3(N__31413),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_9_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_9_12_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_9_12_2  (
            .in0(N__27791),
            .in1(_gnd_net_),
            .in2(N__28758),
            .in3(N__31815),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_9_12_3  (
            .in0(N__32039),
            .in1(N__28483),
            .in2(N__28434),
            .in3(N__28546),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_9_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_9_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_9_12_4  (
            .in0(N__28710),
            .in1(N__27810),
            .in2(_gnd_net_),
            .in3(N__31814),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_12_5 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__28902),
            .in2(N__31128),
            .in3(N__26396),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_9_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_9_12_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_9_12_6  (
            .in0(N__26872),
            .in1(N__27548),
            .in2(_gnd_net_),
            .in3(N__31812),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_9_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_9_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_9_12_7  (
            .in0(N__31813),
            .in1(N__27445),
            .in2(_gnd_net_),
            .in3(N__27980),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_9_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_9_13_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_9_13_1  (
            .in0(N__29604),
            .in1(N__27894),
            .in2(N__29696),
            .in3(N__30464),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_9_13_2  (
            .in0(N__26420),
            .in1(N__26426),
            .in2(N__26381),
            .in3(N__26378),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_9_13_3  (
            .in0(N__26917),
            .in1(N__31748),
            .in2(_gnd_net_),
            .in3(N__29056),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_9_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_9_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_9_13_4  (
            .in0(N__31746),
            .in1(N__31121),
            .in2(_gnd_net_),
            .in3(N__31086),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_9_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_9_13_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_9_13_5  (
            .in0(N__26358),
            .in1(N__31749),
            .in2(_gnd_net_),
            .in3(N__28043),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_9_13_7  (
            .in0(N__29428),
            .in1(N__31747),
            .in2(_gnd_net_),
            .in3(N__29396),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_9_14_0  (
            .in0(N__28233),
            .in1(N__31409),
            .in2(N__28296),
            .in3(N__29055),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_14_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_14_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_9_14_7  (
            .in0(N__28739),
            .in1(N__30767),
            .in2(N__31011),
            .in3(N__28983),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_9_15_0  (
            .in0(N__29252),
            .in1(N__27768),
            .in2(_gnd_net_),
            .in3(N__26414),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__47591),
            .ce(N__29349),
            .sr(N__46886));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_9_15_1  (
            .in0(N__29235),
            .in1(N__27702),
            .in2(_gnd_net_),
            .in3(N__26411),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__47591),
            .ce(N__29349),
            .sr(N__46886));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_9_15_2  (
            .in0(N__29253),
            .in1(N__27627),
            .in2(_gnd_net_),
            .in3(N__26408),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__47591),
            .ce(N__29349),
            .sr(N__46886));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_9_15_3  (
            .in0(N__29236),
            .in1(N__27570),
            .in2(_gnd_net_),
            .in3(N__26405),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__47591),
            .ce(N__29349),
            .sr(N__46886));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_15_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_9_15_4  (
            .in0(N__29254),
            .in1(N__27513),
            .in2(_gnd_net_),
            .in3(N__26402),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__47591),
            .ce(N__29349),
            .sr(N__46886));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_15_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_15_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_9_15_5  (
            .in0(N__29237),
            .in1(N__28206),
            .in2(_gnd_net_),
            .in3(N__26399),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__47591),
            .ce(N__29349),
            .sr(N__46886));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_15_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_15_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_9_15_6  (
            .in0(N__29255),
            .in1(N__28176),
            .in2(_gnd_net_),
            .in3(N__26453),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__47591),
            .ce(N__29349),
            .sr(N__46886));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_15_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_15_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_9_15_7  (
            .in0(N__29238),
            .in1(N__28126),
            .in2(_gnd_net_),
            .in3(N__26450),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__47591),
            .ce(N__29349),
            .sr(N__46886));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_16_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_16_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_9_16_0  (
            .in0(N__29224),
            .in1(N__28071),
            .in2(_gnd_net_),
            .in3(N__26447),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__47585),
            .ce(N__29356),
            .sr(N__46891));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_16_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_16_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_9_16_1  (
            .in0(N__29228),
            .in1(N__28005),
            .in2(_gnd_net_),
            .in3(N__26444),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__47585),
            .ce(N__29356),
            .sr(N__46891));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_16_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_16_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_9_16_2  (
            .in0(N__29221),
            .in1(N__27951),
            .in2(_gnd_net_),
            .in3(N__26441),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__47585),
            .ce(N__29356),
            .sr(N__46891));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_16_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_16_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_9_16_3  (
            .in0(N__29225),
            .in1(N__27925),
            .in2(_gnd_net_),
            .in3(N__26438),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__47585),
            .ce(N__29356),
            .sr(N__46891));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_16_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_16_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_9_16_4  (
            .in0(N__29222),
            .in1(N__27870),
            .in2(_gnd_net_),
            .in3(N__26435),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__47585),
            .ce(N__29356),
            .sr(N__46891));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_16_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_9_16_5  (
            .in0(N__29226),
            .in1(N__28617),
            .in2(_gnd_net_),
            .in3(N__26432),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__47585),
            .ce(N__29356),
            .sr(N__46891));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_16_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_16_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_9_16_6  (
            .in0(N__29223),
            .in1(N__28587),
            .in2(_gnd_net_),
            .in3(N__26429),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__47585),
            .ce(N__29356),
            .sr(N__46891));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_16_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_16_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_9_16_7  (
            .in0(N__29227),
            .in1(N__28521),
            .in2(_gnd_net_),
            .in3(N__26480),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__47585),
            .ce(N__29356),
            .sr(N__46891));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_17_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_17_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_9_17_0  (
            .in0(N__29217),
            .in1(N__28458),
            .in2(_gnd_net_),
            .in3(N__26477),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__47579),
            .ce(N__29348),
            .sr(N__46895));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_17_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_17_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_9_17_1  (
            .in0(N__29248),
            .in1(N__28377),
            .in2(_gnd_net_),
            .in3(N__26474),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__47579),
            .ce(N__29348),
            .sr(N__46895));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_17_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_17_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_9_17_2  (
            .in0(N__29218),
            .in1(N__28350),
            .in2(_gnd_net_),
            .in3(N__26471),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__47579),
            .ce(N__29348),
            .sr(N__46895));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_17_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_9_17_3  (
            .in0(N__29249),
            .in1(N__28323),
            .in2(_gnd_net_),
            .in3(N__26468),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__47579),
            .ce(N__29348),
            .sr(N__46895));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_17_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_17_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_9_17_4  (
            .in0(N__29219),
            .in1(N__28266),
            .in2(_gnd_net_),
            .in3(N__26465),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__47579),
            .ce(N__29348),
            .sr(N__46895));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_17_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_17_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_9_17_5  (
            .in0(N__29250),
            .in1(N__29094),
            .in2(_gnd_net_),
            .in3(N__26462),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__47579),
            .ce(N__29348),
            .sr(N__46895));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_17_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_17_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_9_17_6  (
            .in0(N__29220),
            .in1(N__29025),
            .in2(_gnd_net_),
            .in3(N__26459),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__47579),
            .ce(N__29348),
            .sr(N__46895));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_17_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_17_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_9_17_7  (
            .in0(N__29251),
            .in1(N__28956),
            .in2(_gnd_net_),
            .in3(N__26456),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__47579),
            .ce(N__29348),
            .sr(N__46895));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_18_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_9_18_0  (
            .in0(N__29229),
            .in1(N__28926),
            .in2(_gnd_net_),
            .in3(N__26522),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__47575),
            .ce(N__29357),
            .sr(N__46902));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_18_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_18_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_9_18_1  (
            .in0(N__29233),
            .in1(N__28863),
            .in2(_gnd_net_),
            .in3(N__26519),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__47575),
            .ce(N__29357),
            .sr(N__46902));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_18_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_18_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_9_18_2  (
            .in0(N__29230),
            .in1(N__28839),
            .in2(_gnd_net_),
            .in3(N__26516),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__47575),
            .ce(N__29357),
            .sr(N__46902));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_18_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_9_18_3  (
            .in0(N__29234),
            .in1(N__28782),
            .in2(_gnd_net_),
            .in3(N__26513),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__47575),
            .ce(N__29357),
            .sr(N__46902));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_18_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_18_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_9_18_4  (
            .in0(N__29231),
            .in1(N__28819),
            .in2(_gnd_net_),
            .in3(N__26510),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__47575),
            .ce(N__29357),
            .sr(N__46902));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_18_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_18_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_9_18_5  (
            .in0(N__28798),
            .in1(N__29232),
            .in2(_gnd_net_),
            .in3(N__26507),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47575),
            .ce(N__29357),
            .sr(N__46902));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIPVIS3_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__29299),
            .in2(N__29122),
            .in3(N__29118),
            .lcout(\current_shift_inst.control_input_18 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__33485),
            .in2(_gnd_net_),
            .in3(N__26492),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_19_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__33665),
            .in2(_gnd_net_),
            .in3(N__26483),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_19_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__33647),
            .in2(_gnd_net_),
            .in3(N__26588),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_19_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__33629),
            .in2(_gnd_net_),
            .in3(N__26579),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_19_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__33611),
            .in2(_gnd_net_),
            .in3(N__26570),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_19_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__33593),
            .in2(_gnd_net_),
            .in3(N__26561),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_19_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__33575),
            .in2(_gnd_net_),
            .in3(N__26552),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_20_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__33557),
            .in2(_gnd_net_),
            .in3(N__26543),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_20_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__33833),
            .in2(_gnd_net_),
            .in3(N__26534),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_20_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__33815),
            .in2(_gnd_net_),
            .in3(N__26525),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__34481),
            .in2(_gnd_net_),
            .in3(N__26702),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_20_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__29132),
            .in2(_gnd_net_),
            .in3(N__26693),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_12_c_RNIEEI11_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__37634),
            .in2(_gnd_net_),
            .in3(N__26690),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_9_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_9_20_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26686),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_9_24_0  (
            .in0(_gnd_net_),
            .in1(N__26657),
            .in2(N__26669),
            .in3(N__29557),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__26642),
            .in2(N__26651),
            .in3(N__29535),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_24_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_9_24_2  (
            .in0(N__29514),
            .in1(N__26627),
            .in2(N__26636),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_24_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_9_24_3  (
            .in0(N__29493),
            .in1(N__26612),
            .in2(N__26621),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_24_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_9_24_4  (
            .in0(N__29472),
            .in1(N__26831),
            .in2(N__26606),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_9_24_5  (
            .in0(_gnd_net_),
            .in1(N__26813),
            .in2(N__26825),
            .in3(N__29451),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_24_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_9_24_6  (
            .in0(N__29805),
            .in1(N__26792),
            .in2(N__26807),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_24_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(N__26777),
            .in2(N__26786),
            .in3(N__30623),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_25_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_9_25_0  (
            .in0(N__30642),
            .in1(N__26759),
            .in2(N__26771),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_25_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_9_25_1  (
            .in0(_gnd_net_),
            .in1(N__26744),
            .in2(N__26753),
            .in3(N__30663),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_9_25_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_9_25_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_9_25_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26738),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47556),
            .ce(),
            .sr(N__46930));
    defparam \phase_controller_inst2.S1_LC_9_30_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_30_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_30_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_30_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31178),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47549),
            .ce(),
            .sr(N__46938));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_3_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_3_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_3_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_10_3_5  (
            .in0(N__29734),
            .in1(N__29706),
            .in2(_gnd_net_),
            .in3(N__32007),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_10_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_10_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_10_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_10_4_2  (
            .in0(N__27080),
            .in1(N__28436),
            .in2(_gnd_net_),
            .in3(N__32008),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47689),
            .ce(N__32672),
            .sr(N__46803));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_10_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_10_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_10_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_10_5_4  (
            .in0(N__26847),
            .in1(N__27909),
            .in2(_gnd_net_),
            .in3(N__31983),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47678),
            .ce(N__32648),
            .sr(N__46813));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_10_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_10_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_10_6_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_10_6_0  (
            .in0(N__28160),
            .in1(N__31980),
            .in2(_gnd_net_),
            .in3(N__27023),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__31314),
            .sr(N__46822));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_10_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_10_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_10_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_10_6_1  (
            .in0(N__31975),
            .in1(N__28505),
            .in2(_gnd_net_),
            .in3(N__27005),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__31314),
            .sr(N__46822));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_10_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_10_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_10_6_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_10_6_2  (
            .in0(N__26984),
            .in1(N__31979),
            .in2(_gnd_net_),
            .in3(N__26959),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__31314),
            .sr(N__46822));
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_10_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_10_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_24_LC_10_6_3  (
            .in0(N__31976),
            .in1(N__26921),
            .in2(_gnd_net_),
            .in3(N__29074),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__31314),
            .sr(N__46822));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_10_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_10_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_10_6_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_10_6_4  (
            .in0(N__26896),
            .in1(N__31982),
            .in2(_gnd_net_),
            .in3(N__28570),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__31314),
            .sr(N__46822));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_10_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_10_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_10_6_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_10_6_5  (
            .in0(N__31978),
            .in1(N__27554),
            .in2(_gnd_net_),
            .in3(N__26879),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__31314),
            .sr(N__46822));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_10_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_10_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_10_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_10_6_6  (
            .in0(N__26852),
            .in1(N__27911),
            .in2(_gnd_net_),
            .in3(N__31981),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__31314),
            .sr(N__46822));
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_10_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_10_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_10_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_25_LC_10_6_7  (
            .in0(N__31977),
            .in1(N__27209),
            .in2(_gnd_net_),
            .in3(N__29009),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47669),
            .ce(N__31314),
            .sr(N__46822));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_10_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_10_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__27176),
            .in2(N__27185),
            .in3(N__29838),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_10_7_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_10_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_10_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_10_7_1  (
            .in0(N__29821),
            .in1(N__27170),
            .in2(N__27164),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_10_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_10_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__27155),
            .in2(N__27149),
            .in3(N__30082),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_10_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_10_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(N__27140),
            .in2(N__27131),
            .in3(N__30067),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_10_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_10_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__27119),
            .in2(N__27113),
            .in3(N__30052),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_10_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_10_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(N__27104),
            .in2(N__27098),
            .in3(N__30037),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_10_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_10_7_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_10_7_6  (
            .in0(N__30022),
            .in1(N__31328),
            .in2(N__27089),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_10_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_10_7_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_10_7_7  (
            .in0(N__30007),
            .in1(N__27314),
            .in2(N__29372),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_10_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_10_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__27308),
            .in2(N__27299),
            .in3(N__29993),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_10_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_10_8_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_10_8_1  (
            .in0(N__29974),
            .in1(N__27290),
            .in2(N__27284),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_10_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_10_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__27266),
            .in2(N__27275),
            .in3(N__30244),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_10_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_10_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__27425),
            .in2(N__27260),
            .in3(N__30229),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_10_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_10_8_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_10_8_4  (
            .in0(N__30214),
            .in1(N__30482),
            .in2(N__27251),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_10_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_10_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__27239),
            .in2(N__27230),
            .in3(N__30199),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_10_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_10_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(N__29573),
            .in2(N__27218),
            .in3(N__30184),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_10_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_10_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(N__29633),
            .in2(N__29669),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_10_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_10_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__27359),
            .in2(N__27350),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_10_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_10_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__31520),
            .in2(N__31475),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_10_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_10_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__27335),
            .in2(N__27329),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_10_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_10_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__27455),
            .in2(N__27491),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_10_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_10_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__27416),
            .in2(N__27410),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_10_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_10_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__27368),
            .in2(N__27842),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_10_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_10_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_LUT4_0_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__29870),
            .in2(N__29945),
            .in3(N__27317),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27494),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_10_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_10_10_0  (
            .in0(N__30334),
            .in1(N__27482),
            .in2(N__27470),
            .in3(N__30315),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_10_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_10_10_1  (
            .in0(N__27481),
            .in1(N__27469),
            .in2(N__30317),
            .in3(N__30333),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_10_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_10_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_10_10_4  (
            .in0(N__27449),
            .in1(N__27982),
            .in2(_gnd_net_),
            .in3(N__31905),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47622),
            .ce(N__31310),
            .sr(N__46849));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_10_7 .LUT_INIT=16'b1000111010101111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_10_10_7  (
            .in0(N__27379),
            .in1(N__30497),
            .in2(N__30274),
            .in3(N__30295),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_10_11_0  (
            .in0(N__30493),
            .in1(N__27380),
            .in2(N__30275),
            .in3(N__30294),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_10_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_10_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_10_11_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_27_LC_10_11_1  (
            .in0(N__28901),
            .in1(N__31774),
            .in2(_gnd_net_),
            .in3(N__27398),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47612),
            .ce(N__31308),
            .sr(N__46855));
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_10_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_10_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_28_LC_10_11_2  (
            .in0(N__31772),
            .in1(N__31132),
            .in2(_gnd_net_),
            .in3(N__31096),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47612),
            .ce(N__31308),
            .sr(N__46855));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_11_3 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_10_11_3  (
            .in0(N__27850),
            .in1(N__30571),
            .in2(N__30596),
            .in3(N__27826),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_11_4 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_10_11_4  (
            .in0(N__30591),
            .in1(N__30570),
            .in2(N__27830),
            .in3(N__27851),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_10_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_10_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_10_11_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_29_LC_10_11_5  (
            .in0(N__31023),
            .in1(N__31775),
            .in2(_gnd_net_),
            .in3(N__31046),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47612),
            .ce(N__31308),
            .sr(N__46855));
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_10_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_10_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_10_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_31_LC_10_11_6  (
            .in0(N__31773),
            .in1(N__28717),
            .in2(_gnd_net_),
            .in3(N__27818),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47612),
            .ce(N__31308),
            .sr(N__46855));
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_10_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_30_LC_10_11_7  (
            .in0(N__28759),
            .in1(N__27790),
            .in2(_gnd_net_),
            .in3(N__31776),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47612),
            .ce(N__31308),
            .sr(N__46855));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_12_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__27773),
            .in2(N__27632),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47601),
            .ce(N__28684),
            .sr(N__46861));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__27571),
            .in2(N__27710),
            .in3(N__27635),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47601),
            .ce(N__28684),
            .sr(N__46861));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__27631),
            .in2(N__27520),
            .in3(N__27575),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47601),
            .ce(N__28684),
            .sr(N__46861));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__27572),
            .in2(N__28213),
            .in3(N__27524),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47601),
            .ce(N__28684),
            .sr(N__46861));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__28183),
            .in2(N__27521),
            .in3(N__27497),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47601),
            .ce(N__28684),
            .sr(N__46861));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(N__28132),
            .in2(N__28214),
            .in3(N__28190),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47601),
            .ce(N__28684),
            .sr(N__46861));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(N__28078),
            .in2(N__28187),
            .in3(N__28136),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47601),
            .ce(N__28684),
            .sr(N__46861));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(N__28133),
            .in2(N__28018),
            .in3(N__28085),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47601),
            .ce(N__28684),
            .sr(N__46861));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__27952),
            .in2(N__28082),
            .in3(N__28022),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47593),
            .ce(N__28685),
            .sr(N__46866));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__27931),
            .in2(N__28019),
            .in3(N__27956),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47593),
            .ce(N__28685),
            .sr(N__46866));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__27953),
            .in2(N__27877),
            .in3(N__27935),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47593),
            .ce(N__28685),
            .sr(N__46866));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(N__27932),
            .in2(N__28624),
            .in3(N__27881),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47593),
            .ce(N__28685),
            .sr(N__46866));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(N__28594),
            .in2(N__27878),
            .in3(N__27854),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47593),
            .ce(N__28685),
            .sr(N__46866));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_13_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(N__28528),
            .in2(N__28625),
            .in3(N__28601),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47593),
            .ce(N__28685),
            .sr(N__46866));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_13_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_13_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(N__28465),
            .in2(N__28598),
            .in3(N__28535),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47593),
            .ce(N__28685),
            .sr(N__46866));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_13_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__28384),
            .in2(N__28532),
            .in3(N__28472),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47593),
            .ce(N__28685),
            .sr(N__46866));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_14_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_14_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__28351),
            .in2(N__28469),
            .in3(N__28388),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47586),
            .ce(N__28676),
            .sr(N__46870));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_14_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_14_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__28385),
            .in2(N__28330),
            .in3(N__28355),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47586),
            .ce(N__28676),
            .sr(N__46870));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_14_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_14_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__28352),
            .in2(N__28273),
            .in3(N__28334),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47586),
            .ce(N__28676),
            .sr(N__46870));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_14_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_14_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__29095),
            .in2(N__28331),
            .in3(N__28277),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47586),
            .ce(N__28676),
            .sr(N__46870));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_14_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_14_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__29032),
            .in2(N__28274),
            .in3(N__28217),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47586),
            .ce(N__28676),
            .sr(N__46870));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_14_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_14_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(N__28963),
            .in2(N__29099),
            .in3(N__29039),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47586),
            .ce(N__28676),
            .sr(N__46870));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_14_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_14_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__28933),
            .in2(N__29036),
            .in3(N__28970),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47586),
            .ce(N__28676),
            .sr(N__46870));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_14_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_14_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__28871),
            .in2(N__28967),
            .in3(N__28940),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47586),
            .ce(N__28676),
            .sr(N__46870));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_15_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_15_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__28840),
            .in2(N__28937),
            .in3(N__28874),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47580),
            .ce(N__28675),
            .sr(N__46874));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_15_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_15_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__28870),
            .in2(N__28783),
            .in3(N__28844),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47580),
            .ce(N__28675),
            .sr(N__46874));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_15_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_15_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__28841),
            .in2(N__28823),
            .in3(N__28805),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47580),
            .ce(N__28675),
            .sr(N__46874));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_15_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_15_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__28802),
            .in2(N__28784),
            .in3(N__28724),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47580),
            .ce(N__28675),
            .sr(N__46874));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_15_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28721),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47580),
            .ce(N__28675),
            .sr(N__46874));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_10_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_10_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_10_16_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_10_16_4  (
            .in0(N__29432),
            .in1(N__29407),
            .in2(_gnd_net_),
            .in3(N__32003),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47577),
            .ce(N__31307),
            .sr(N__46880));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_17_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_17_0 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_10_17_0  (
            .in0(N__30915),
            .in1(N__29279),
            .in2(_gnd_net_),
            .in3(N__32959),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_203_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_17_1.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_17_1.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MAX_D2_LC_10_17_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MAX_D2_LC_10_17_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29318),
            .lcout(il_max_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47570),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_17_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_10_17_2  (
            .in0(N__34331),
            .in1(N__32729),
            .in2(_gnd_net_),
            .in3(N__37589),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_10_17_3  (
            .in0(N__29278),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_10_18_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_10_18_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_10_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30719),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30677),
            .ce(),
            .sr(N__46892));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_19_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_10_19_2  (
            .in0(N__37632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37631),
            .lcout(\current_shift_inst.N_1304_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_10_23_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_10_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__29515),
            .in2(_gnd_net_),
            .in3(N__29556),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_10_23_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_10_23_5 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_10_23_5  (
            .in0(N__29473),
            .in1(N__29494),
            .in2(N__29564),
            .in3(N__29536),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_10_23_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_10_23_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_10_23_6  (
            .in0(N__30602),
            .in1(N__29807),
            .in2(N__29561),
            .in3(N__29453),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_10_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_10_24_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_10_24_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_10_24_0  (
            .in0(N__29775),
            .in1(N__29558),
            .in2(_gnd_net_),
            .in3(N__29540),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_10_24_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__47555),
            .ce(),
            .sr(N__46918));
    defparam \pwm_generator_inst.counter_1_LC_10_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_10_24_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_10_24_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_10_24_1  (
            .in0(N__29771),
            .in1(N__29537),
            .in2(_gnd_net_),
            .in3(N__29519),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__47555),
            .ce(),
            .sr(N__46918));
    defparam \pwm_generator_inst.counter_2_LC_10_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_10_24_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_10_24_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_10_24_2  (
            .in0(N__29776),
            .in1(N__29516),
            .in2(_gnd_net_),
            .in3(N__29498),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__47555),
            .ce(),
            .sr(N__46918));
    defparam \pwm_generator_inst.counter_3_LC_10_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_10_24_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_10_24_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_10_24_3  (
            .in0(N__29772),
            .in1(N__29495),
            .in2(_gnd_net_),
            .in3(N__29477),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__47555),
            .ce(),
            .sr(N__46918));
    defparam \pwm_generator_inst.counter_4_LC_10_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_10_24_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_10_24_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_10_24_4  (
            .in0(N__29777),
            .in1(N__29474),
            .in2(_gnd_net_),
            .in3(N__29456),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__47555),
            .ce(),
            .sr(N__46918));
    defparam \pwm_generator_inst.counter_5_LC_10_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_10_24_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_10_24_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_10_24_5  (
            .in0(N__29773),
            .in1(N__29452),
            .in2(_gnd_net_),
            .in3(N__29435),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__47555),
            .ce(),
            .sr(N__46918));
    defparam \pwm_generator_inst.counter_6_LC_10_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_10_24_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_10_24_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_10_24_6  (
            .in0(N__29778),
            .in1(N__29806),
            .in2(_gnd_net_),
            .in3(N__29789),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__47555),
            .ce(),
            .sr(N__46918));
    defparam \pwm_generator_inst.counter_7_LC_10_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_10_24_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_10_24_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_10_24_7  (
            .in0(N__29774),
            .in1(N__30622),
            .in2(_gnd_net_),
            .in3(N__29786),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__47555),
            .ce(),
            .sr(N__46918));
    defparam \pwm_generator_inst.counter_8_LC_10_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_10_25_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_10_25_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_10_25_0  (
            .in0(N__29780),
            .in1(N__30643),
            .in2(_gnd_net_),
            .in3(N__29783),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_10_25_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__47552),
            .ce(),
            .sr(N__46922));
    defparam \pwm_generator_inst.counter_9_LC_10_25_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_10_25_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_10_25_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_10_25_1  (
            .in0(N__30664),
            .in1(N__29779),
            .in2(_gnd_net_),
            .in3(N__29738),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47552),
            .ce(),
            .sr(N__46922));
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_4_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_4_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_RNO_0_LC_11_4_5  (
            .in0(N__31203),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31173),
            .lcout(\phase_controller_inst2.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_11_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_11_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_11_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_11_5_2  (
            .in0(N__29735),
            .in1(N__29714),
            .in2(_gnd_net_),
            .in3(N__32005),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47670),
            .ce(N__31316),
            .sr(N__46804));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_6_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_11_6_0  (
            .in0(N__30139),
            .in1(N__29645),
            .in2(N__30170),
            .in3(N__29654),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_6_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_11_6_1  (
            .in0(N__29653),
            .in1(N__30169),
            .in2(N__30143),
            .in3(N__29644),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_11_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_11_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_11_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_11_6_6  (
            .in0(N__29624),
            .in1(N__29588),
            .in2(_gnd_net_),
            .in3(N__32004),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47656),
            .ce(N__31315),
            .sr(N__46814));
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_7_0 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_RNISIH31_30_LC_11_7_0  (
            .in0(N__30550),
            .in1(N__30524),
            .in2(N__29924),
            .in3(N__29889),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_hc.un4_running_df30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_7_1 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIEABO2_28_LC_11_7_1  (
            .in0(N__29935),
            .in1(N__32230),
            .in2(N__29960),
            .in3(N__29957),
            .lcout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_7_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29948),
            .in3(N__32295),
            .lcout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_7_3 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_RNISIH31_0_30_LC_11_7_3  (
            .in0(N__29919),
            .in1(N__30519),
            .in2(N__29893),
            .in3(N__30549),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3_28_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__32296),
            .in2(_gnd_net_),
            .in3(N__29860),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI6OQI3Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_7_5 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_11_7_5  (
            .in0(N__29920),
            .in1(N__30520),
            .in2(N__29894),
            .in3(N__30551),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_7_6 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_11_7_6  (
            .in0(N__32172),
            .in1(N__29861),
            .in2(N__29846),
            .in3(N__32297),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47646),
            .ce(),
            .sr(N__46823));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__29852),
            .in2(N__29845),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_11_8_1  (
            .in0(N__32177),
            .in1(N__29822),
            .in2(_gnd_net_),
            .in3(N__29810),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__47634),
            .ce(),
            .sr(N__46829));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_8_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_11_8_2  (
            .in0(N__32181),
            .in1(N__30083),
            .in2(N__30092),
            .in3(N__30071),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__47634),
            .ce(),
            .sr(N__46829));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_11_8_3  (
            .in0(N__32178),
            .in1(N__30068),
            .in2(_gnd_net_),
            .in3(N__30056),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__47634),
            .ce(),
            .sr(N__46829));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_11_8_4  (
            .in0(N__32182),
            .in1(N__30053),
            .in2(_gnd_net_),
            .in3(N__30041),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__47634),
            .ce(),
            .sr(N__46829));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_11_8_5  (
            .in0(N__32179),
            .in1(N__30038),
            .in2(_gnd_net_),
            .in3(N__30026),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__47634),
            .ce(),
            .sr(N__46829));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_11_8_6  (
            .in0(N__32183),
            .in1(N__30023),
            .in2(_gnd_net_),
            .in3(N__30011),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__47634),
            .ce(),
            .sr(N__46829));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_11_8_7  (
            .in0(N__32180),
            .in1(N__30008),
            .in2(_gnd_net_),
            .in3(N__29996),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__47634),
            .ce(),
            .sr(N__46829));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_11_9_0  (
            .in0(N__32176),
            .in1(N__29992),
            .in2(_gnd_net_),
            .in3(N__29978),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__47623),
            .ce(),
            .sr(N__46837));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_11_9_1  (
            .in0(N__32188),
            .in1(N__29975),
            .in2(_gnd_net_),
            .in3(N__29963),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__47623),
            .ce(),
            .sr(N__46837));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_11_9_2  (
            .in0(N__32173),
            .in1(N__30245),
            .in2(_gnd_net_),
            .in3(N__30233),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__47623),
            .ce(),
            .sr(N__46837));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_11_9_3  (
            .in0(N__32189),
            .in1(N__30230),
            .in2(_gnd_net_),
            .in3(N__30218),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__47623),
            .ce(),
            .sr(N__46837));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_11_9_4  (
            .in0(N__32174),
            .in1(N__30215),
            .in2(_gnd_net_),
            .in3(N__30203),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__47623),
            .ce(),
            .sr(N__46837));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_11_9_5  (
            .in0(N__32190),
            .in1(N__30200),
            .in2(_gnd_net_),
            .in3(N__30188),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__47623),
            .ce(),
            .sr(N__46837));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_11_9_6  (
            .in0(N__32175),
            .in1(N__30185),
            .in2(_gnd_net_),
            .in3(N__30173),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__47623),
            .ce(),
            .sr(N__46837));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_11_9_7  (
            .in0(N__32191),
            .in1(N__30160),
            .in2(_gnd_net_),
            .in3(N__30146),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__47623),
            .ce(),
            .sr(N__46837));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_11_10_0  (
            .in0(N__32184),
            .in1(N__30138),
            .in2(_gnd_net_),
            .in3(N__30119),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__47613),
            .ce(),
            .sr(N__46844));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_11_10_1  (
            .in0(N__32165),
            .in1(N__30109),
            .in2(_gnd_net_),
            .in3(N__30095),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__47613),
            .ce(),
            .sr(N__46844));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_11_10_2  (
            .in0(N__32185),
            .in1(N__30409),
            .in2(_gnd_net_),
            .in3(N__30395),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__47613),
            .ce(),
            .sr(N__46844));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_11_10_3  (
            .in0(N__32166),
            .in1(N__31510),
            .in2(_gnd_net_),
            .in3(N__30392),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__47613),
            .ce(),
            .sr(N__46844));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_11_10_4  (
            .in0(N__32186),
            .in1(N__31492),
            .in2(_gnd_net_),
            .in3(N__30389),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__47613),
            .ce(),
            .sr(N__46844));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_11_10_5  (
            .in0(N__32167),
            .in1(N__30376),
            .in2(_gnd_net_),
            .in3(N__30362),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__47613),
            .ce(),
            .sr(N__46844));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_11_10_6  (
            .in0(N__32187),
            .in1(N__30352),
            .in2(_gnd_net_),
            .in3(N__30338),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__47613),
            .ce(),
            .sr(N__46844));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_11_10_7  (
            .in0(N__32168),
            .in1(N__30335),
            .in2(_gnd_net_),
            .in3(N__30320),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__47613),
            .ce(),
            .sr(N__46844));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_11_11_0  (
            .in0(N__32109),
            .in1(N__30316),
            .in2(_gnd_net_),
            .in3(N__30299),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__47602),
            .ce(),
            .sr(N__46850));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_11_11_1  (
            .in0(N__32113),
            .in1(N__30296),
            .in2(_gnd_net_),
            .in3(N__30278),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__47602),
            .ce(),
            .sr(N__46850));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_11_11_2  (
            .in0(N__32110),
            .in1(N__30270),
            .in2(_gnd_net_),
            .in3(N__30248),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__47602),
            .ce(),
            .sr(N__46850));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_11_11_3  (
            .in0(N__32114),
            .in1(N__30595),
            .in2(_gnd_net_),
            .in3(N__30575),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__47602),
            .ce(),
            .sr(N__46850));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_11_11_4  (
            .in0(N__32111),
            .in1(N__30572),
            .in2(_gnd_net_),
            .in3(N__30554),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__47602),
            .ce(),
            .sr(N__46850));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_11_11_5  (
            .in0(N__32115),
            .in1(N__30548),
            .in2(_gnd_net_),
            .in3(N__30530),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__47602),
            .ce(),
            .sr(N__46850));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_11_11_6  (
            .in0(N__32112),
            .in1(N__30518),
            .in2(_gnd_net_),
            .in3(N__30527),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47602),
            .ce(),
            .sr(N__46850));
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_11_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_11_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_26_LC_11_12_6  (
            .in0(N__31833),
            .in1(N__30745),
            .in2(_gnd_net_),
            .in3(N__30775),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47594),
            .ce(N__31309),
            .sr(N__46856));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_11_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_11_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_11_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_11_12_7  (
            .in0(N__30435),
            .in1(N__30466),
            .in2(_gnd_net_),
            .in3(N__31834),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47594),
            .ce(N__31309),
            .sr(N__46856));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_11_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_11_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_11_13_4  (
            .in0(N__30439),
            .in1(N__30465),
            .in2(_gnd_net_),
            .in3(N__31943),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_11_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_11_14_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNO_LC_11_14_1  (
            .in0(N__44192),
            .in1(N__39281),
            .in2(N__45051),
            .in3(N__42190),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_11_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_11_14_4 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNO_LC_11_14_4  (
            .in0(N__42799),
            .in1(N__45003),
            .in2(N__39374),
            .in3(N__44193),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_11_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_ns_i_a2_1_LC_11_15_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_ns_i_a2_1_LC_11_15_1  (
            .in0(N__30810),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34662),
            .lcout(state_ns_i_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_15_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_15_4 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__33444),
            .in2(N__30725),
            .in3(N__30694),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_205_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_15_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_15_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_11_15_5  (
            .in0(N__30768),
            .in1(N__30744),
            .in2(_gnd_net_),
            .in3(N__31937),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_15_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_15_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__33443),
            .in2(_gnd_net_),
            .in3(N__30693),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_204_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_11_16_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_11_16_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_11_16_5 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_11_16_5  (
            .in0(N__33445),
            .in1(N__30724),
            .in2(_gnd_net_),
            .in3(N__30695),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47571),
            .ce(),
            .sr(N__46875));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_17_1 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_11_17_1  (
            .in0(N__45035),
            .in1(N__40022),
            .in2(N__44416),
            .in3(N__43441),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_17_6 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_11_17_6  (
            .in0(N__44355),
            .in1(N__40072),
            .in2(N__43309),
            .in3(N__45036),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_18_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_18_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30720),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__30676),
            .ce(),
            .sr(N__46887));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_11_23_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_11_23_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_11_23_7  (
            .in0(N__30665),
            .in1(N__30644),
            .in2(_gnd_net_),
            .in3(N__30618),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_24_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_24_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_11_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32947),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32926),
            .ce(),
            .sr(N__46914));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_6.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_11_30_6 (
            .in0(N__30887),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_12_3_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNIG7JF_2_LC_12_3_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst2.state_RNIG7JF_2_LC_12_3_1  (
            .in0(N__30862),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31275),
            .lcout(\phase_controller_inst2.state_RNIG7JFZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_12_3_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_12_3_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_12_3_3  (
            .in0(N__30861),
            .in1(N__31276),
            .in2(N__33010),
            .in3(N__31238),
            .lcout(\phase_controller_inst2.start_timer_tr_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_LC_12_4_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_12_4_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_12_4_3 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_12_4_3  (
            .in0(N__30869),
            .in1(N__32891),
            .in2(N__32878),
            .in3(N__34689),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47668),
            .ce(),
            .sr(N__46792));
    defparam \phase_controller_inst2.state_2_LC_12_4_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_12_4_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_12_4_5 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \phase_controller_inst2.state_2_LC_12_4_5  (
            .in0(N__31204),
            .in1(N__31169),
            .in2(N__31280),
            .in3(N__30863),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47668),
            .ce(),
            .sr(N__46792));
    defparam \phase_controller_inst2.start_timer_hc_LC_12_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_12_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_12_4_6 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_12_4_6  (
            .in0(N__34688),
            .in1(N__30838),
            .in2(N__32261),
            .in3(N__30848),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47668),
            .ce(),
            .sr(N__46792));
    defparam \phase_controller_inst2.state_1_LC_12_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_12_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_12_5_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \phase_controller_inst2.state_1_LC_12_5_3  (
            .in0(N__31237),
            .in1(N__33003),
            .in2(_gnd_net_),
            .in3(N__30842),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47655),
            .ce(),
            .sr(N__46797));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_12_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32879),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47655),
            .ce(),
            .sr(N__46797));
    defparam \phase_controller_inst2.state_0_LC_12_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_12_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_12_5_7 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \phase_controller_inst2.state_0_LC_12_5_7  (
            .in0(N__31236),
            .in1(N__33002),
            .in2(N__32852),
            .in3(N__32903),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47655),
            .ce(),
            .sr(N__46797));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_6_2 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_6_2  (
            .in0(N__33077),
            .in1(N__33050),
            .in2(N__34728),
            .in3(N__34092),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47645),
            .ce(),
            .sr(N__46805));
    defparam \phase_controller_inst2.state_3_LC_12_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_12_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_12_6_5 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \phase_controller_inst2.state_3_LC_12_6_5  (
            .in0(N__31208),
            .in1(N__32890),
            .in2(N__31174),
            .in3(N__33791),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47645),
            .ce(),
            .sr(N__46805));
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_12_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_12_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_12_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_28_LC_12_7_5  (
            .in0(N__31133),
            .in1(N__31097),
            .in2(_gnd_net_),
            .in3(N__32006),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47633),
            .ce(N__32656),
            .sr(N__46815));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_8_0 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_8_0  (
            .in0(N__30992),
            .in1(N__30982),
            .in2(N__30964),
            .in3(N__30941),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_8_2  (
            .in0(N__31024),
            .in1(N__31984),
            .in2(_gnd_net_),
            .in3(N__31039),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_12_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_12_8_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_29_LC_12_8_3  (
            .in0(N__31986),
            .in1(_gnd_net_),
            .in2(N__31028),
            .in3(N__31025),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47621),
            .ce(N__32594),
            .sr(N__46824));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_12_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_12_8_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_12_8_4  (
            .in0(N__30991),
            .in1(N__30983),
            .in2(N__30965),
            .in3(N__30940),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_12_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_12_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_12_8_5  (
            .in0(N__31985),
            .in1(N__31371),
            .in2(_gnd_net_),
            .in3(N__31339),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_12_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_12_8_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_12_8_6  (
            .in0(N__31372),
            .in1(_gnd_net_),
            .in2(N__31535),
            .in3(N__31987),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47621),
            .ce(N__32594),
            .sr(N__46824));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_9_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_12_9_0  (
            .in0(N__31382),
            .in1(N__31463),
            .in2(N__31511),
            .in3(N__31491),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_9_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_12_9_1  (
            .in0(N__31462),
            .in1(N__31509),
            .in2(N__31493),
            .in3(N__31381),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_12_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_12_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_20_LC_12_9_2  (
            .in0(N__32045),
            .in1(N__31561),
            .in2(_gnd_net_),
            .in3(N__31958),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47611),
            .ce(N__31313),
            .sr(N__46830));
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_12_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_12_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_21_LC_12_9_3  (
            .in0(N__31956),
            .in1(N__31454),
            .in2(_gnd_net_),
            .in3(N__31424),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47611),
            .ce(N__31313),
            .sr(N__46830));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_12_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_12_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_12_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_12_9_7  (
            .in0(N__31957),
            .in1(N__31373),
            .in2(_gnd_net_),
            .in3(N__31340),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47611),
            .ce(N__31313),
            .sr(N__46830));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_2 .LUT_INIT=16'b1101110000001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_12_10_2  (
            .in0(N__31252),
            .in1(N__31274),
            .in2(N__32294),
            .in3(N__32229),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47600),
            .ce(),
            .sr(N__46838));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_12_10_3  (
            .in0(N__32266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47600),
            .ce(),
            .sr(N__46838));
    defparam \phase_controller_inst2.stoper_hc.running_LC_12_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_12_10_5 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_12_10_5  (
            .in0(N__32228),
            .in1(N__31253),
            .in2(N__32312),
            .in3(N__32286),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47600),
            .ce(),
            .sr(N__46838));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_11_1 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_12_11_1  (
            .in0(N__42040),
            .in1(N__42062),
            .in2(N__38674),
            .in3(N__47191),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47592),
            .ce(),
            .sr(N__46845));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_11_2 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_12_11_2  (
            .in0(N__32497),
            .in1(N__32399),
            .in2(N__32384),
            .in3(N__32328),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47592),
            .ce(),
            .sr(N__46845));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_11_4 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_12_11_4  (
            .in0(N__32221),
            .in1(N__32308),
            .in2(_gnd_net_),
            .in3(N__32262),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_12_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_12_12_5  (
            .in0(N__32267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32231),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_12_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_12_12_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_12_12_7  (
            .in0(N__31560),
            .in1(N__32041),
            .in2(_gnd_net_),
            .in3(N__31938),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42261),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_13_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__44191),
            .in2(N__31538),
            .in3(N__33199),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42416),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47576),
            .ce(N__43572),
            .sr(N__46862));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_14_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_12_14_4  (
            .in0(N__44189),
            .in1(N__44919),
            .in2(N__39326),
            .in3(N__42226),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_14_5 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_12_14_5  (
            .in0(N__42227),
            .in1(N__39325),
            .in2(N__45029),
            .in3(N__44190),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__34262),
            .in2(N__33464),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__45157),
            .in2(N__45131),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__44858),
            .in2(N__32693),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__32684),
            .in2(N__45004),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__44862),
            .in2(N__36359),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__36098),
            .in2(N__45005),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__44866),
            .in2(N__39770),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__32678),
            .in2(N__45006),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__44870),
            .in2(N__36068),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__33275),
            .in2(N__45007),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__44874),
            .in2(N__33290),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__33296),
            .in2(N__45008),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__44878),
            .in2(N__33269),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__33545),
            .in2(N__45009),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__44882),
            .in2(N__33539),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__33281),
            .in2(N__45010),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__44886),
            .in2(N__33515),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__40205),
            .in2(N__45011),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__44890),
            .in2(N__33530),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__33521),
            .in2(N__45012),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(N__44894),
            .in2(N__33506),
            .in3(N__32720),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(N__40214),
            .in2(N__45013),
            .in3(N__32717),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_12_17_6  (
            .in0(_gnd_net_),
            .in1(N__44898),
            .in2(N__32714),
            .in3(N__32702),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(N__33497),
            .in2(N__45014),
            .in3(N__32699),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(N__45015),
            .in2(N__33803),
            .in3(N__32696),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(N__32783),
            .in2(N__45052),
            .in3(N__32777),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__45019),
            .in2(N__34439),
            .in3(N__32774),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(N__36470),
            .in2(N__45053),
            .in3(N__32771),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(N__45023),
            .in2(N__40232),
            .in3(N__32768),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__33677),
            .in2(N__45054),
            .in3(N__32765),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__45027),
            .in2(N__45113),
            .in3(N__32762),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_18_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_12_18_7  (
            .in0(N__45028),
            .in1(N__44391),
            .in2(_gnd_net_),
            .in3(N__32759),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_20_0.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_20_0.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D2_LC_12_20_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 SB_DFF_inst_PH1_MIN_D2_LC_12_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32735),
            .lcout(il_min_comp1_D2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47560),
            .ce(),
            .sr(_gnd_net_));
    defparam SB_DFF_inst_PH1_MIN_D1_LC_12_20_5.C_ON=1'b0;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_12_20_5.SEQ_MODE=4'b1000;
    defparam SB_DFF_inst_PH1_MIN_D1_LC_12_20_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 SB_DFF_inst_PH1_MIN_D1_LC_12_20_5 (
            .in0(N__32756),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(il_min_comp1_D1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47560),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.S2_LC_12_21_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_12_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33011),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47557),
            .ce(),
            .sr(N__46896));
    defparam \delay_measurement_inst.start_timer_hc_LC_12_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_12_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32946),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32927),
            .ce(),
            .sr(N__46909));
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1 .C_ON=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1 .SEQ_MODE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_RNO_LC_12_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46958),
            .lcout(\pll_inst.red_c_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_13_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNI9M3O_0_LC_13_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.state_RNI9M3O_0_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(N__32847),
            .in2(_gnd_net_),
            .in3(N__32902),
            .lcout(\phase_controller_inst2.state_RNI9M3OZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_5_6 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_13_5_6  (
            .in0(N__32801),
            .in1(N__32830),
            .in2(_gnd_net_),
            .in3(N__32870),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_5_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_5_7  (
            .in0(N__32871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32802),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_3 .LUT_INIT=16'b1101000011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_13_6_3  (
            .in0(N__35296),
            .in1(N__32851),
            .in2(N__32813),
            .in3(N__33076),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47657),
            .ce(),
            .sr(N__46798));
    defparam \phase_controller_inst2.stoper_tr.running_LC_13_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_13_7_3 .LUT_INIT=16'b1101010111110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_13_7_3  (
            .in0(N__32812),
            .in1(N__35297),
            .in2(N__32831),
            .in3(N__33079),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47647),
            .ce(),
            .sr(N__46806));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_7_4 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNISIOB3_28_LC_13_7_4  (
            .in0(N__35332),
            .in1(N__32811),
            .in2(N__33038),
            .in3(N__35315),
            .lcout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33083),
            .in3(N__33078),
            .lcout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_8_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_8_1  (
            .in0(N__41524),
            .in1(N__41503),
            .in2(_gnd_net_),
            .in3(N__48116),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34_28_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__33080),
            .in2(_gnd_net_),
            .in3(N__33049),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI5PG34Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_13_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_13_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_13_8_4  (
            .in0(N__48117),
            .in1(N__37216),
            .in2(_gnd_net_),
            .in3(N__37260),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_9_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_0_30_LC_13_9_0  (
            .in0(N__34206),
            .in1(N__34023),
            .in2(N__33119),
            .in3(N__33025),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_9_1 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_RNI8K5A1_30_LC_13_9_1  (
            .in0(N__33024),
            .in1(N__34207),
            .in2(N__34030),
            .in3(N__33114),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_df30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_13_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_13_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_30_LC_13_9_2  (
            .in0(N__41063),
            .in1(N__48187),
            .in2(_gnd_net_),
            .in3(N__34001),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47624),
            .ce(N__45954),
            .sr(N__46825));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_9_3 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_13_9_3  (
            .in0(N__33026),
            .in1(N__34208),
            .in2(N__34031),
            .in3(N__33118),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_13_9_4  (
            .in0(N__34273),
            .in1(N__48186),
            .in2(_gnd_net_),
            .in3(N__38457),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_13_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_13_9_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_13_9_5  (
            .in0(N__48189),
            .in1(_gnd_net_),
            .in2(N__33014),
            .in3(N__38458),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47624),
            .ce(N__45954),
            .sr(N__46825));
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_13_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_13_9_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_31_LC_13_9_6  (
            .in0(N__34295),
            .in1(N__48188),
            .in2(_gnd_net_),
            .in3(N__38356),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47624),
            .ce(N__45954),
            .sr(N__46825));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_13_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_13_9_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_13_9_7  (
            .in0(N__41504),
            .in1(N__41520),
            .in2(N__48206),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47624),
            .ce(N__45954),
            .sr(N__46825));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_13_10_0  (
            .in0(N__33405),
            .in1(N__35604),
            .in2(_gnd_net_),
            .in3(N__33104),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__47614),
            .ce(N__33245),
            .sr(N__46831));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_13_10_1  (
            .in0(N__33397),
            .in1(N__35577),
            .in2(_gnd_net_),
            .in3(N__33101),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__47614),
            .ce(N__33245),
            .sr(N__46831));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_13_10_2  (
            .in0(N__33406),
            .in1(N__35547),
            .in2(_gnd_net_),
            .in3(N__33098),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__47614),
            .ce(N__33245),
            .sr(N__46831));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_13_10_3  (
            .in0(N__33398),
            .in1(N__35526),
            .in2(_gnd_net_),
            .in3(N__33095),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__47614),
            .ce(N__33245),
            .sr(N__46831));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_13_10_4  (
            .in0(N__33407),
            .in1(N__35502),
            .in2(_gnd_net_),
            .in3(N__33092),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__47614),
            .ce(N__33245),
            .sr(N__46831));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_13_10_5  (
            .in0(N__33399),
            .in1(N__35472),
            .in2(_gnd_net_),
            .in3(N__33089),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__47614),
            .ce(N__33245),
            .sr(N__46831));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_13_10_6  (
            .in0(N__33408),
            .in1(N__35453),
            .in2(_gnd_net_),
            .in3(N__33086),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__47614),
            .ce(N__33245),
            .sr(N__46831));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_13_10_7  (
            .in0(N__33400),
            .in1(N__35427),
            .in2(_gnd_net_),
            .in3(N__33146),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__47614),
            .ce(N__33245),
            .sr(N__46831));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_13_11_0  (
            .in0(N__33396),
            .in1(N__35394),
            .in2(_gnd_net_),
            .in3(N__33143),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__47603),
            .ce(N__33244),
            .sr(N__46839));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_13_11_1  (
            .in0(N__33404),
            .in1(N__35823),
            .in2(_gnd_net_),
            .in3(N__33140),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__47603),
            .ce(N__33244),
            .sr(N__46839));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_13_11_2  (
            .in0(N__33393),
            .in1(N__35793),
            .in2(_gnd_net_),
            .in3(N__33137),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__47603),
            .ce(N__33244),
            .sr(N__46839));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_13_11_3  (
            .in0(N__33401),
            .in1(N__35769),
            .in2(_gnd_net_),
            .in3(N__33134),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__47603),
            .ce(N__33244),
            .sr(N__46839));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_13_11_4  (
            .in0(N__33394),
            .in1(N__35739),
            .in2(_gnd_net_),
            .in3(N__33131),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__47603),
            .ce(N__33244),
            .sr(N__46839));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_13_11_5  (
            .in0(N__33402),
            .in1(N__35715),
            .in2(_gnd_net_),
            .in3(N__33128),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__47603),
            .ce(N__33244),
            .sr(N__46839));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_13_11_6  (
            .in0(N__33395),
            .in1(N__35688),
            .in2(_gnd_net_),
            .in3(N__33125),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__47603),
            .ce(N__33244),
            .sr(N__46839));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_13_11_7  (
            .in0(N__33403),
            .in1(N__35666),
            .in2(_gnd_net_),
            .in3(N__33122),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__47603),
            .ce(N__33244),
            .sr(N__46839));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_13_12_0  (
            .in0(N__33415),
            .in1(N__35637),
            .in2(_gnd_net_),
            .in3(N__33173),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__47595),
            .ce(N__33237),
            .sr(N__46846));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_13_12_1  (
            .in0(N__33419),
            .in1(N__36030),
            .in2(_gnd_net_),
            .in3(N__33170),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__47595),
            .ce(N__33237),
            .sr(N__46846));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_13_12_2  (
            .in0(N__33416),
            .in1(N__36001),
            .in2(_gnd_net_),
            .in3(N__33167),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__47595),
            .ce(N__33237),
            .sr(N__46846));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_13_12_3  (
            .in0(N__33420),
            .in1(N__35976),
            .in2(_gnd_net_),
            .in3(N__33164),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__47595),
            .ce(N__33237),
            .sr(N__46846));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_13_12_4  (
            .in0(N__33417),
            .in1(N__35955),
            .in2(_gnd_net_),
            .in3(N__33161),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__47595),
            .ce(N__33237),
            .sr(N__46846));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_13_12_5  (
            .in0(N__33421),
            .in1(N__35931),
            .in2(_gnd_net_),
            .in3(N__33158),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__47595),
            .ce(N__33237),
            .sr(N__46846));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_13_12_6  (
            .in0(N__33418),
            .in1(N__35901),
            .in2(_gnd_net_),
            .in3(N__33155),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__47595),
            .ce(N__33237),
            .sr(N__46846));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_13_12_7  (
            .in0(N__33422),
            .in1(N__35874),
            .in2(_gnd_net_),
            .in3(N__33152),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__47595),
            .ce(N__33237),
            .sr(N__46846));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_13_13_0  (
            .in0(N__33409),
            .in1(N__35844),
            .in2(_gnd_net_),
            .in3(N__33149),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__47587),
            .ce(N__33236),
            .sr(N__46851));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_13_13_1  (
            .in0(N__33413),
            .in1(N__36279),
            .in2(_gnd_net_),
            .in3(N__33260),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__47587),
            .ce(N__33236),
            .sr(N__46851));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_13_13_2  (
            .in0(N__33410),
            .in1(N__36235),
            .in2(_gnd_net_),
            .in3(N__33257),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__47587),
            .ce(N__33236),
            .sr(N__46851));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_13_13_3  (
            .in0(N__33414),
            .in1(N__36192),
            .in2(_gnd_net_),
            .in3(N__33254),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__47587),
            .ce(N__33236),
            .sr(N__46851));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_13_13_4  (
            .in0(N__33411),
            .in1(N__36253),
            .in2(_gnd_net_),
            .in3(N__33251),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__47587),
            .ce(N__33236),
            .sr(N__46851));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_13_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_13_13_5  (
            .in0(N__36211),
            .in1(N__33412),
            .in2(_gnd_net_),
            .in3(N__33248),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47587),
            .ce(N__33236),
            .sr(N__46851));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40154),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47581),
            .ce(N__43571),
            .sr(N__46857));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33194),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_2 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_14_2  (
            .in0(N__33195),
            .in1(_gnd_net_),
            .in2(N__33203),
            .in3(N__42383),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42415),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47581),
            .ce(N__43571),
            .sr(N__46857));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_14_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__44239),
            .in2(N__33200),
            .in3(N__33179),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_13_14_6  (
            .in0(N__37501),
            .in1(N__37759),
            .in2(_gnd_net_),
            .in3(N__33473),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_13_14_7  (
            .in0(N__37760),
            .in1(_gnd_net_),
            .in2(N__33467),
            .in3(N__33463),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_15_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNO_LC_13_15_0  (
            .in0(N__44925),
            .in1(N__44200),
            .in2(N__39710),
            .in3(N__43183),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_15_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33449),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_15_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNO_LC_13_15_2  (
            .in0(N__44924),
            .in1(N__44196),
            .in2(N__39620),
            .in3(N__42631),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_15_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNO_LC_13_15_3  (
            .in0(N__44195),
            .in1(N__44923),
            .in2(N__42671),
            .in3(N__39664),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_15_4 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNO_LC_13_15_4  (
            .in0(N__43070),
            .in1(N__44199),
            .in2(N__45030),
            .in3(N__39571),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_15_5 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNO_LC_13_15_5  (
            .in0(N__44194),
            .in1(N__39493),
            .in2(N__42719),
            .in3(N__44931),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_15_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNO_LC_13_15_6  (
            .in0(N__44926),
            .in1(N__44197),
            .in2(N__39709),
            .in3(N__43184),
            .lcout(\current_shift_inst.un38_control_input_cry_12_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_15_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNO_LC_13_15_7  (
            .in0(N__44198),
            .in1(N__44927),
            .in2(N__39757),
            .in3(N__43147),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNO_LC_13_16_0  (
            .in0(N__44291),
            .in1(N__44935),
            .in2(N__43121),
            .in3(N__44061),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_1 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_13_16_1  (
            .in0(N__44932),
            .in1(N__40018),
            .in2(N__43442),
            .in3(N__44297),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_16_2 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNO_LC_13_16_2  (
            .in0(N__44293),
            .in1(N__42956),
            .in2(N__39925),
            .in3(N__44937),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_16_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNO_LC_13_16_3  (
            .in0(N__44938),
            .in1(N__44294),
            .in2(N__43907),
            .in3(N__42931),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_16_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNO_LC_13_16_4  (
            .in0(N__44292),
            .in1(N__44936),
            .in2(N__40121),
            .in3(N__43031),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_13_16_6 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_13_16_6  (
            .in0(N__44295),
            .in1(N__39878),
            .in2(N__43520),
            .in3(N__44934),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_16_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_13_16_7  (
            .in0(N__44933),
            .in1(N__44296),
            .in2(N__43397),
            .in3(N__39971),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_17_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_13_17_0  (
            .in0(N__33491),
            .in1(N__34316),
            .in2(_gnd_net_),
            .in3(N__37593),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_17_1 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_13_17_1  (
            .in0(N__44948),
            .in1(N__44012),
            .in2(N__43727),
            .in3(N__44298),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_17_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_13_17_2  (
            .in0(N__33671),
            .in1(N__34415),
            .in2(_gnd_net_),
            .in3(N__37594),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_17_3 .LUT_INIT=16'b0101000001011111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_13_17_3  (
            .in0(N__34403),
            .in1(_gnd_net_),
            .in2(N__37621),
            .in3(N__33653),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_17_4 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_13_17_4  (
            .in0(N__33635),
            .in1(N__34391),
            .in2(_gnd_net_),
            .in3(N__37598),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_17_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_13_17_5  (
            .in0(N__37599),
            .in1(N__33617),
            .in2(_gnd_net_),
            .in3(N__34382),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_17_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_13_17_6  (
            .in0(N__33599),
            .in1(N__34373),
            .in2(_gnd_net_),
            .in3(N__37600),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_17_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_13_17_7  (
            .in0(N__37601),
            .in1(N__34364),
            .in2(_gnd_net_),
            .in3(N__33581),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_13_18_0  (
            .in0(N__33563),
            .in1(N__34355),
            .in2(_gnd_net_),
            .in3(N__37622),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_18_1 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_13_18_1  (
            .in0(N__34343),
            .in1(N__37624),
            .in2(_gnd_net_),
            .in3(N__33839),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_18_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_13_18_2  (
            .in0(N__33821),
            .in1(N__34508),
            .in2(_gnd_net_),
            .in3(N__37623),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_18_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_13_18_7  (
            .in0(N__44417),
            .in1(N__40348),
            .in2(N__45046),
            .in3(N__43355),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_13_19_1 .LUT_INIT=16'b1101000011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_13_19_1  (
            .in0(N__42145),
            .in1(N__38079),
            .in2(N__45506),
            .in3(N__42044),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47562),
            .ce(),
            .sr(N__46881));
    defparam \phase_controller_inst1.state_3_LC_13_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_13_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_13_19_3 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \phase_controller_inst1.state_3_LC_13_19_3  (
            .in0(N__36693),
            .in1(N__38020),
            .in2(N__33716),
            .in3(N__33787),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47562),
            .ce(),
            .sr(N__46881));
    defparam \phase_controller_inst1.start_timer_hc_LC_13_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_19_7 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_13_19_7  (
            .in0(N__33722),
            .in1(N__34637),
            .in2(N__34691),
            .in3(N__33741),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47562),
            .ce(),
            .sr(N__46881));
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_20_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_RNO_0_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__36678),
            .in2(_gnd_net_),
            .in3(N__33708),
            .lcout(\phase_controller_inst1.start_timer_hc_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_2_LC_13_22_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_13_22_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_13_22_6 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \phase_controller_inst1.state_2_LC_13_22_6  (
            .in0(N__33715),
            .in1(N__36636),
            .in2(N__34619),
            .in3(N__36696),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47558),
            .ce(),
            .sr(N__46897));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__34529),
            .in2(_gnd_net_),
            .in3(N__34843),
            .lcout(\current_shift_inst.timer_s1.N_162_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_LC_13_24_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_13_24_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_13_24_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_13_24_3  (
            .in0(N__34895),
            .in1(N__34534),
            .in2(_gnd_net_),
            .in3(N__34842),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47553),
            .ce(),
            .sr(N__46905));
    defparam \phase_controller_inst1.S1_LC_13_25_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_13_25_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_13_25_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_13_25_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36695),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47551),
            .ce(),
            .sr(N__46910));
    defparam \current_shift_inst.start_timer_s1_LC_13_25_7 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_13_25_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_13_25_7 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_13_25_7  (
            .in0(N__34860),
            .in1(N__34893),
            .in2(_gnd_net_),
            .in3(N__36694),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47551),
            .ce(),
            .sr(N__46910));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_14_6_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_14_6_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_14_6_0  (
            .in0(N__38160),
            .in1(N__38213),
            .in2(N__37262),
            .in3(N__37280),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35615),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47671),
            .ce(N__36167),
            .sr(N__46793));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_6_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35588),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47671),
            .ce(N__36167),
            .sr(N__46793));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_14_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_14_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_14_6_4  (
            .in0(N__37309),
            .in1(N__37281),
            .in2(_gnd_net_),
            .in3(N__48144),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_7_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_14_7_0  (
            .in0(N__33979),
            .in1(N__33955),
            .in2(N__33893),
            .in3(N__33848),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_7_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_14_7_1  (
            .in0(N__33847),
            .in1(N__33980),
            .in2(N__33959),
            .in3(N__33889),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_14_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_14_7_2  (
            .in0(N__42599),
            .in1(N__48184),
            .in2(_gnd_net_),
            .in3(N__41855),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47658),
            .ce(N__45952),
            .sr(N__46799));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_14_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_14_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_14_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_14_7_3  (
            .in0(N__48181),
            .in1(N__41936),
            .in2(_gnd_net_),
            .in3(N__41904),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47658),
            .ce(N__45952),
            .sr(N__46799));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_14_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_14_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_14_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_14_7_4  (
            .in0(N__37261),
            .in1(N__48185),
            .in2(_gnd_net_),
            .in3(N__37212),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47658),
            .ce(N__45952),
            .sr(N__46799));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_14_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_14_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_14_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_14_7_5  (
            .in0(N__48182),
            .in1(N__38265),
            .in2(_gnd_net_),
            .in3(N__36896),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47658),
            .ce(N__45952),
            .sr(N__46799));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_14_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_14_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_14_7_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_14_7_7  (
            .in0(N__48183),
            .in1(N__38762),
            .in2(_gnd_net_),
            .in3(N__38798),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47658),
            .ce(N__45952),
            .sr(N__46799));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__33881),
            .in2(N__34733),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_14_8_1  (
            .in0(N__34145),
            .in1(N__35072),
            .in2(_gnd_net_),
            .in3(N__33875),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__47648),
            .ce(),
            .sr(N__46807));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_8_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_14_8_2  (
            .in0(N__34142),
            .in1(N__35045),
            .in2(N__33872),
            .in3(N__33860),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__47648),
            .ce(),
            .sr(N__46807));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_14_8_3  (
            .in0(N__34146),
            .in1(N__35015),
            .in2(_gnd_net_),
            .in3(N__33857),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__47648),
            .ce(),
            .sr(N__46807));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_14_8_4  (
            .in0(N__34143),
            .in1(N__34988),
            .in2(_gnd_net_),
            .in3(N__33854),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__47648),
            .ce(),
            .sr(N__46807));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_14_8_5  (
            .in0(N__34147),
            .in1(N__34964),
            .in2(_gnd_net_),
            .in3(N__33851),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__47648),
            .ce(),
            .sr(N__46807));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_14_8_6  (
            .in0(N__34144),
            .in1(N__34937),
            .in2(_gnd_net_),
            .in3(N__33920),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__47648),
            .ce(),
            .sr(N__46807));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_14_8_7  (
            .in0(N__34148),
            .in1(N__34916),
            .in2(_gnd_net_),
            .in3(N__33917),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__47648),
            .ce(),
            .sr(N__46807));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_14_9_0  (
            .in0(N__34179),
            .in1(N__35273),
            .in2(_gnd_net_),
            .in3(N__33914),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__47635),
            .ce(),
            .sr(N__46816));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_14_9_1  (
            .in0(N__34181),
            .in1(N__35252),
            .in2(_gnd_net_),
            .in3(N__33911),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__47635),
            .ce(),
            .sr(N__46816));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_14_9_2  (
            .in0(N__34176),
            .in1(N__35231),
            .in2(_gnd_net_),
            .in3(N__33908),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__47635),
            .ce(),
            .sr(N__46816));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_14_9_3  (
            .in0(N__34182),
            .in1(N__35213),
            .in2(_gnd_net_),
            .in3(N__33905),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__47635),
            .ce(),
            .sr(N__46816));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_14_9_4  (
            .in0(N__34177),
            .in1(N__35182),
            .in2(_gnd_net_),
            .in3(N__33902),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__47635),
            .ce(),
            .sr(N__46816));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_14_9_5  (
            .in0(N__34183),
            .in1(N__35144),
            .in2(_gnd_net_),
            .in3(N__33899),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__47635),
            .ce(),
            .sr(N__46816));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_14_9_6  (
            .in0(N__34178),
            .in1(N__35114),
            .in2(_gnd_net_),
            .in3(N__33896),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__47635),
            .ce(),
            .sr(N__46816));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_14_9_7  (
            .in0(N__34184),
            .in1(N__34767),
            .in2(_gnd_net_),
            .in3(N__33986),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__47635),
            .ce(),
            .sr(N__46816));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_14_10_0  (
            .in0(N__34161),
            .in1(N__34795),
            .in2(_gnd_net_),
            .in3(N__33983),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__47625),
            .ce(),
            .sr(N__46826));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_14_10_1  (
            .in0(N__34165),
            .in1(N__33978),
            .in2(_gnd_net_),
            .in3(N__33962),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__47625),
            .ce(),
            .sr(N__46826));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_14_10_2  (
            .in0(N__34162),
            .in1(N__33954),
            .in2(_gnd_net_),
            .in3(N__33938),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__47625),
            .ce(),
            .sr(N__46826));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_14_10_3  (
            .in0(N__34166),
            .in1(N__36829),
            .in2(_gnd_net_),
            .in3(N__33935),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__47625),
            .ce(),
            .sr(N__46826));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_14_10_4  (
            .in0(N__34163),
            .in1(N__36801),
            .in2(_gnd_net_),
            .in3(N__33932),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__47625),
            .ce(),
            .sr(N__46826));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_14_10_5  (
            .in0(N__34167),
            .in1(N__36946),
            .in2(_gnd_net_),
            .in3(N__33929),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__47625),
            .ce(),
            .sr(N__46826));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_14_10_6  (
            .in0(N__34164),
            .in1(N__36970),
            .in2(_gnd_net_),
            .in3(N__33926),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__47625),
            .ce(),
            .sr(N__46826));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_14_10_7  (
            .in0(N__34168),
            .in1(N__45406),
            .in2(_gnd_net_),
            .in3(N__33923),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__47625),
            .ce(),
            .sr(N__46826));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_14_11_0  (
            .in0(N__34169),
            .in1(N__45436),
            .in2(_gnd_net_),
            .in3(N__34223),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__47615),
            .ce(),
            .sr(N__46832));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_14_11_1  (
            .in0(N__34173),
            .in1(N__45361),
            .in2(_gnd_net_),
            .in3(N__34220),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__47615),
            .ce(),
            .sr(N__46832));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_14_11_2  (
            .in0(N__34170),
            .in1(N__45337),
            .in2(_gnd_net_),
            .in3(N__34217),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__47615),
            .ce(),
            .sr(N__46832));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_14_11_3  (
            .in0(N__34174),
            .in1(N__45243),
            .in2(_gnd_net_),
            .in3(N__34214),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__47615),
            .ce(),
            .sr(N__46832));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_14_11_4  (
            .in0(N__34171),
            .in1(N__45276),
            .in2(_gnd_net_),
            .in3(N__34211),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__47615),
            .ce(),
            .sr(N__46832));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_14_11_5  (
            .in0(N__34175),
            .in1(N__34205),
            .in2(_gnd_net_),
            .in3(N__34187),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__47615),
            .ce(),
            .sr(N__46832));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_14_11_6  (
            .in0(N__34172),
            .in1(N__34015),
            .in2(_gnd_net_),
            .in3(N__34034),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47615),
            .ce(),
            .sr(N__46832));
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_14_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_14_12_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_0_30_LC_14_12_0  (
            .in0(N__39525),
            .in1(N__38841),
            .in2(N__39170),
            .in3(N__38817),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_14_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_14_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_14_12_1  (
            .in0(N__41045),
            .in1(N__33997),
            .in2(_gnd_net_),
            .in3(N__48194),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_14_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_14_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_14_12_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_30_LC_14_12_2  (
            .in0(N__48195),
            .in1(_gnd_net_),
            .in2(N__34298),
            .in3(N__41046),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47604),
            .ce(N__47208),
            .sr(N__46840));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_14_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_14_12_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_14_12_3  (
            .in0(N__38342),
            .in1(N__34291),
            .in2(_gnd_net_),
            .in3(N__48193),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(elapsed_time_ns_1_RNI0CQBB_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_14_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_14_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_14_12_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_31_LC_14_12_4  (
            .in0(N__48196),
            .in1(_gnd_net_),
            .in2(N__34280),
            .in3(N__38343),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47604),
            .ce(N__47208),
            .sr(N__46840));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_14_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_14_12_5 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_14_12_5  (
            .in0(N__38842),
            .in1(N__39169),
            .in2(N__38824),
            .in3(N__39526),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_14_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_14_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_14_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_14_12_7  (
            .in0(N__34277),
            .in1(N__48197),
            .in2(_gnd_net_),
            .in3(N__38444),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47604),
            .ce(N__47208),
            .sr(N__46840));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__34261),
            .in2(N__34250),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__45150),
            .in2(N__43610),
            .in3(N__45071),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2  (
            .in0(N__45072),
            .in1(N__44552),
            .in2(N__34238),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__34460),
            .in2(N__44775),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_LC_14_13_4  (
            .in0(_gnd_net_),
            .in1(N__44556),
            .in2(N__36086),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__36074),
            .in2(N__44776),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_13_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_LC_14_13_6  (
            .in0(_gnd_net_),
            .in1(N__44560),
            .in2(N__43628),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_13_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(N__36320),
            .in2(N__44777),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__44564),
            .in2(N__36311),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__36344),
            .in2(N__44778),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__44568),
            .in2(N__36437),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__36053),
            .in2(N__44779),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__44572),
            .in2(N__34307),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__36302),
            .in2(N__44780),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__44576),
            .in2(N__36335),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__36326),
            .in2(N__44781),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__44782),
            .in2(N__36296),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__34451),
            .in2(N__44969),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__44786),
            .in2(N__36410),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__36428),
            .in2(N__44970),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__44790),
            .in2(N__36422),
            .in3(N__34319),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__42428),
            .in2(N__44971),
            .in3(N__34427),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__44794),
            .in2(N__34424),
            .in3(N__34406),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__36392),
            .in2(N__44972),
            .in3(N__34394),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__44798),
            .in2(N__36386),
            .in3(N__34385),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__36458),
            .in2(N__44973),
            .in3(N__34376),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__44802),
            .in2(N__36401),
            .in3(N__34367),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__36365),
            .in2(N__44974),
            .in3(N__34358),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__44806),
            .in2(N__36374),
            .in3(N__34346),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__34466),
            .in2(N__44975),
            .in3(N__34334),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__44810),
            .in2(N__44078),
            .in3(N__34499),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7  (
            .in0(N__42479),
            .in1(N__34496),
            .in2(N__37633),
            .in3(N__34484),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39434),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39474),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_14_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_14_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_14_17_4  (
            .in0(N__44400),
            .in1(N__44008),
            .in2(N__45043),
            .in3(N__43726),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_17_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNO_LC_14_17_6  (
            .in0(N__44398),
            .in1(N__39273),
            .in2(N__45044),
            .in3(N__42191),
            .lcout(\current_shift_inst.un38_control_input_cry_3_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_17_7 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNO_LC_14_17_7  (
            .in0(N__42998),
            .in1(N__44979),
            .in2(N__43967),
            .in3(N__44399),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_3  (
            .in0(N__40191),
            .in1(N__44407),
            .in2(N__45045),
            .in3(N__43262),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39596),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40052),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39642),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_LC_14_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_14_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_14_20_1 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_14_20_1  (
            .in0(N__34690),
            .in1(N__34544),
            .in2(N__45539),
            .in3(N__38024),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47563),
            .ce(),
            .sr(N__46882));
    defparam \phase_controller_inst1.state_0_LC_14_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_14_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_14_20_5 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \phase_controller_inst1.state_0_LC_14_20_5  (
            .in0(N__38046),
            .in1(N__38080),
            .in2(N__34574),
            .in3(N__36576),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47563),
            .ce(),
            .sr(N__46882));
    defparam \phase_controller_inst1.state_1_LC_14_20_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_14_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_14_20_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst1.state_1_LC_14_20_6  (
            .in0(N__36577),
            .in1(N__34572),
            .in2(_gnd_net_),
            .in3(N__34633),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47563),
            .ce(),
            .sr(N__46882));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_14_22_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_14_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNIE87F_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(N__36634),
            .in2(_gnd_net_),
            .in3(N__34614),
            .lcout(\phase_controller_inst1.time_passed_RNIE87F ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_22_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34535),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_23_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_23_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_14_23_1  (
            .in0(N__36635),
            .in1(N__34615),
            .in2(N__34573),
            .in3(N__36578),
            .lcout(\phase_controller_inst1.start_timer_tr_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_24_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_14_24_1  (
            .in0(N__34892),
            .in1(N__34533),
            .in2(_gnd_net_),
            .in3(N__34838),
            .lcout(\current_shift_inst.timer_s1.N_163_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.stop_timer_s1_LC_14_25_1 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_14_25_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_14_25_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_14_25_1  (
            .in0(N__34894),
            .in1(N__36703),
            .in2(N__34844),
            .in3(N__34861),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47554),
            .ce(),
            .sr(N__46906));
    defparam \phase_controller_inst1.S2_LC_14_27_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_14_27_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_14_27_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.S2_LC_14_27_5  (
            .in0(N__36587),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47550),
            .ce(),
            .sr(N__46915));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_5_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_15_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_15_5_0  (
            .in0(N__38120),
            .in1(N__38159),
            .in2(_gnd_net_),
            .in3(N__48180),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47690),
            .ce(N__47219),
            .sr(N__46785));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_6_0 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_15_6_0  (
            .in0(N__34750),
            .in1(N__36863),
            .in2(N__34780),
            .in3(N__34802),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_6_1 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_15_6_1  (
            .in0(N__34801),
            .in1(N__34751),
            .in2(N__34781),
            .in3(N__36862),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_15_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_15_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_15_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_15_6_2  (
            .in0(N__41454),
            .in1(N__41420),
            .in2(_gnd_net_),
            .in3(N__48147),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47679),
            .ce(N__45953),
            .sr(N__46788));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_15_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_15_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_15_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_15_6_4  (
            .in0(N__42518),
            .in1(N__42545),
            .in2(_gnd_net_),
            .in3(N__48146),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47679),
            .ce(N__45953),
            .sr(N__46788));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_15_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_15_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_15_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_15_6_5  (
            .in0(N__48145),
            .in1(N__37305),
            .in2(_gnd_net_),
            .in3(N__37282),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47679),
            .ce(N__45953),
            .sr(N__46788));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_15_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_15_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_15_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_15_6_6  (
            .in0(N__38191),
            .in1(N__38217),
            .in2(_gnd_net_),
            .in3(N__48148),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47679),
            .ce(N__45953),
            .sr(N__46788));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_15_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_15_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(N__34742),
            .in2(N__34700),
            .in3(N__34729),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_15_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_15_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_15_7_1  (
            .in0(N__35071),
            .in1(N__35060),
            .in2(N__35054),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_15_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_15_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__36875),
            .in2(N__35033),
            .in3(N__35044),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_15_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_15_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(N__35024),
            .in2(N__35003),
            .in3(N__35014),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_15_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_15_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(N__34994),
            .in2(N__34976),
            .in3(N__34987),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_15_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_15_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__36869),
            .in2(N__34952),
            .in3(N__34963),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_15_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_15_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__34943),
            .in2(N__34925),
            .in3(N__34936),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_15_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_15_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__37007),
            .in2(N__34904),
            .in3(N__34915),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_15_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_15_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__35261),
            .in2(N__37001),
            .in3(N__35272),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_15_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_15_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__36992),
            .in2(N__35240),
            .in3(N__35251),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_15_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_15_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__35219),
            .in2(N__36905),
            .in3(N__35230),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_15_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_15_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__35201),
            .in2(N__37106),
            .in3(N__35212),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_15_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_15_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__35195),
            .in2(N__35168),
            .in3(N__35183),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_15_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_15_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__35159),
            .in2(N__35132),
            .in3(N__35143),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_15_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_15_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(N__35123),
            .in2(N__35102),
            .in3(N__35113),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_15_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_15_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__35093),
            .in2(N__35084),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_15_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_15_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(N__35369),
            .in2(N__35360),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_15_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_15_9_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__36773),
            .in2(N__36851),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_15_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_15_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__36932),
            .in2(N__36986),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_15_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_15_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__45392),
            .in2(N__43781),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_15_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_15_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__45380),
            .in2(N__45323),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_15_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_15_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__45302),
            .in2(N__45731),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_15_9_6  (
            .in0(_gnd_net_),
            .in1(N__35345),
            .in2(N__35336),
            .in3(N__35303),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35300),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__35611),
            .in2(N__35554),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47636),
            .ce(N__36166),
            .sr(N__46817));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__35527),
            .in2(N__35587),
            .in3(N__35558),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47636),
            .ce(N__36166),
            .sr(N__46817));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__35503),
            .in2(N__35555),
            .in3(N__35531),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47636),
            .ce(N__36166),
            .sr(N__46817));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__35528),
            .in2(N__35479),
            .in3(N__35510),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47636),
            .ce(N__36166),
            .sr(N__46817));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__35451),
            .in2(N__35507),
            .in3(N__35483),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47636),
            .ce(N__36166),
            .sr(N__46817));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__35428),
            .in2(N__35480),
            .in3(N__35456),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47636),
            .ce(N__36166),
            .sr(N__46817));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__35452),
            .in2(N__35405),
            .in3(N__35435),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47636),
            .ce(N__36166),
            .sr(N__46817));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__35824),
            .in2(N__35432),
            .in3(N__35408),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47636),
            .ce(N__36166),
            .sr(N__46817));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__35794),
            .in2(N__35404),
            .in3(N__35372),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47626),
            .ce(N__36158),
            .sr(N__46827));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__35770),
            .in2(N__35825),
            .in3(N__35798),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47626),
            .ce(N__36158),
            .sr(N__46827));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__35795),
            .in2(N__35746),
            .in3(N__35777),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47626),
            .ce(N__36158),
            .sr(N__46827));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__35716),
            .in2(N__35774),
            .in3(N__35750),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47626),
            .ce(N__36158),
            .sr(N__46827));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__35689),
            .in2(N__35747),
            .in3(N__35723),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47626),
            .ce(N__36158),
            .sr(N__46827));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__35664),
            .in2(N__35720),
            .in3(N__35696),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47626),
            .ce(N__36158),
            .sr(N__46827));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(N__35644),
            .in2(N__35693),
            .in3(N__35669),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47626),
            .ce(N__36158),
            .sr(N__46827));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__35665),
            .in2(N__36041),
            .in3(N__35648),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47626),
            .ce(N__36158),
            .sr(N__46827));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__36000),
            .in2(N__35645),
            .in3(N__35618),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47616),
            .ce(N__36159),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__35977),
            .in2(N__36040),
            .in3(N__36008),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47616),
            .ce(N__36159),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__35956),
            .in2(N__36005),
            .in3(N__35981),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47616),
            .ce(N__36159),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__35978),
            .in2(N__35936),
            .in3(N__35960),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47616),
            .ce(N__36159),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__35957),
            .in2(N__35908),
            .in3(N__35939),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47616),
            .ce(N__36159),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__35935),
            .in2(N__35881),
            .in3(N__35912),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47616),
            .ce(N__36159),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(N__35851),
            .in2(N__35909),
            .in3(N__35885),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47616),
            .ce(N__36159),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__36286),
            .in2(N__35882),
            .in3(N__35858),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47616),
            .ce(N__36159),
            .sr(N__46833));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__36234),
            .in2(N__35855),
            .in3(N__35828),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47605),
            .ce(N__36157),
            .sr(N__46841));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__36193),
            .in2(N__36287),
            .in3(N__36257),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47605),
            .ce(N__36157),
            .sr(N__46841));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__36254),
            .in2(N__36239),
            .in3(N__36215),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47605),
            .ce(N__36157),
            .sr(N__46841));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__36212),
            .in2(N__36197),
            .in3(N__36173),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47605),
            .ce(N__36157),
            .sr(N__46841));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36170),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47605),
            .ce(N__36157),
            .sr(N__46841));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_14_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNO_LC_15_14_0  (
            .in0(N__44625),
            .in1(N__44278),
            .in2(N__39823),
            .in3(N__42845),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_14_1 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNO_LC_15_14_1  (
            .in0(N__44280),
            .in1(N__39407),
            .in2(N__42890),
            .in3(N__44623),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_14_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNO_LC_15_14_2  (
            .in0(N__44624),
            .in1(N__44281),
            .in2(N__39824),
            .in3(N__42844),
            .lcout(\current_shift_inst.un38_control_input_cry_5_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_14_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNO_LC_15_14_3  (
            .in0(N__44279),
            .in1(N__44626),
            .in2(N__42760),
            .in3(N__39447),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_4 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNO_LC_15_14_4  (
            .in0(N__44622),
            .in1(N__44282),
            .in2(N__39619),
            .in3(N__42632),
            .lcout(\current_shift_inst.un38_control_input_cry_11_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_14_6 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNO_LC_15_14_6  (
            .in0(N__39406),
            .in1(N__44277),
            .in2(N__42889),
            .in3(N__44627),
            .lcout(\current_shift_inst.un38_control_input_cry_4_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_14_7 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_14_7  (
            .in0(N__45194),
            .in1(N__45211),
            .in2(_gnd_net_),
            .in3(N__42380),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_15_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNO_LC_15_15_0  (
            .in0(N__44361),
            .in1(N__39489),
            .in2(N__44996),
            .in3(N__42715),
            .lcout(\current_shift_inst.un38_control_input_cry_9_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_15_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNO_LC_15_15_1  (
            .in0(N__44063),
            .in1(N__44364),
            .in2(N__43117),
            .in3(N__44829),
            .lcout(\current_shift_inst.un38_control_input_cry_14_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_15_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNO_LC_15_15_2  (
            .in0(N__44365),
            .in1(N__43069),
            .in2(N__44994),
            .in3(N__39567),
            .lcout(\current_shift_inst.un38_control_input_cry_15_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_15_3 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNO_LC_15_15_3  (
            .in0(N__42803),
            .in1(N__44834),
            .in2(N__39373),
            .in3(N__44359),
            .lcout(\current_shift_inst.un38_control_input_cry_7_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_15_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNO_LC_15_15_4  (
            .in0(N__44360),
            .in1(N__39448),
            .in2(N__44995),
            .in3(N__42761),
            .lcout(\current_shift_inst.un38_control_input_cry_8_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_15_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_15_15_5 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNO_LC_15_15_5  (
            .in0(N__43151),
            .in1(N__44828),
            .in2(N__39758),
            .in3(N__44363),
            .lcout(\current_shift_inst.un38_control_input_cry_13_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_15_6 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNO_LC_15_15_6  (
            .in0(N__44833),
            .in1(N__43027),
            .in2(N__44419),
            .in3(N__40120),
            .lcout(\current_shift_inst.un38_control_input_cry_16_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_15_7 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNO_LC_15_15_7  (
            .in0(N__42670),
            .in1(N__44827),
            .in2(N__39665),
            .in3(N__44362),
            .lcout(\current_shift_inst.un38_control_input_cry_10_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_16_0 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNO_LC_15_16_0  (
            .in0(N__44852),
            .in1(N__43900),
            .in2(N__42932),
            .in3(N__44402),
            .lcout(\current_shift_inst.un38_control_input_cry_19_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_15_16_1  (
            .in0(N__44403),
            .in1(N__39876),
            .in2(N__44998),
            .in3(N__43516),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_16_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNO_LC_15_16_2  (
            .in0(N__44851),
            .in1(N__44401),
            .in2(N__39926),
            .in3(N__42955),
            .lcout(\current_shift_inst.un38_control_input_cry_18_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_16_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_16_3  (
            .in0(N__44406),
            .in1(N__40192),
            .in2(N__44999),
            .in3(N__43261),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_16_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_15_16_4  (
            .in0(N__42381),
            .in1(N__42927),
            .in2(_gnd_net_),
            .in3(N__43899),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_16_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_16_5  (
            .in0(N__44404),
            .in1(N__39970),
            .in2(N__44997),
            .in3(N__43396),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_16_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_15_16_6  (
            .in0(N__44850),
            .in1(N__44405),
            .in2(N__40352),
            .in3(N__43348),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_17_0 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_15_17_0  (
            .in0(N__44389),
            .in1(N__45033),
            .in2(N__43754),
            .in3(N__40260),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_17_1 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_17_1  (
            .in0(N__45031),
            .in1(N__40303),
            .in2(N__44429),
            .in3(N__43216),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_17_3 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_15_17_3  (
            .in0(N__45032),
            .in1(N__40304),
            .in2(N__44428),
            .in3(N__43217),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39350),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_6 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_6  (
            .in0(N__44388),
            .in1(N__40065),
            .in2(N__43310),
            .in3(N__45034),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_18_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__40567),
            .in2(N__40153),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__47572),
            .ce(N__43570),
            .sr(N__46867));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__43595),
            .in2(N__40547),
            .in3(N__36452),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__47572),
            .ce(N__43570),
            .sr(N__46867));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__40568),
            .in2(N__40516),
            .in3(N__36449),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__47572),
            .ce(N__43570),
            .sr(N__46867));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__40546),
            .in2(N__40489),
            .in3(N__36446),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__47572),
            .ce(N__43570),
            .sr(N__46867));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__40462),
            .in2(N__40517),
            .in3(N__36443),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__47572),
            .ce(N__43570),
            .sr(N__46867));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__40441),
            .in2(N__40490),
            .in3(N__36440),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__47572),
            .ce(N__43570),
            .sr(N__46867));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__40463),
            .in2(N__40420),
            .in3(N__36497),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__47572),
            .ce(N__43570),
            .sr(N__46867));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__40442),
            .in2(N__40387),
            .in3(N__36494),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__47572),
            .ce(N__43570),
            .sr(N__46867));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__40783),
            .in2(N__40421),
            .in3(N__36491),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__47567),
            .ce(N__43569),
            .sr(N__46871));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__40762),
            .in2(N__40388),
            .in3(N__36488),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__47567),
            .ce(N__43569),
            .sr(N__46871));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__40784),
            .in2(N__40742),
            .in3(N__36485),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__47567),
            .ce(N__43569),
            .sr(N__46871));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__40763),
            .in2(N__40715),
            .in3(N__36482),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__47567),
            .ce(N__43569),
            .sr(N__46871));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__40741),
            .in2(N__40687),
            .in3(N__36479),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__47567),
            .ce(N__43569),
            .sr(N__46871));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__40714),
            .in2(N__40660),
            .in3(N__36476),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__47567),
            .ce(N__43569),
            .sr(N__46871));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__40633),
            .in2(N__40688),
            .in3(N__36473),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__47567),
            .ce(N__43569),
            .sr(N__46871));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__40600),
            .in2(N__40661),
            .in3(N__36524),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__47567),
            .ce(N__43569),
            .sr(N__46871));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(N__41017),
            .in2(N__40634),
            .in3(N__36521),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__47565),
            .ce(N__43568),
            .sr(N__46876));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__40993),
            .in2(N__40601),
            .in3(N__36518),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__47565),
            .ce(N__43568),
            .sr(N__46876));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(N__41018),
            .in2(N__40969),
            .in3(N__36515),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__47565),
            .ce(N__43568),
            .sr(N__46876));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__40942),
            .in2(N__40997),
            .in3(N__36512),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__47565),
            .ce(N__43568),
            .sr(N__46876));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_15_20_4  (
            .in0(_gnd_net_),
            .in1(N__40921),
            .in2(N__40970),
            .in3(N__36509),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__47565),
            .ce(N__43568),
            .sr(N__46876));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(N__40943),
            .in2(N__40900),
            .in3(N__36506),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__47565),
            .ce(N__43568),
            .sr(N__46876));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__40922),
            .in2(N__40874),
            .in3(N__36503),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__47565),
            .ce(N__43568),
            .sr(N__46876));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_15_20_7  (
            .in0(_gnd_net_),
            .in1(N__40837),
            .in2(N__40901),
            .in3(N__36500),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__47565),
            .ce(N__43568),
            .sr(N__46876));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_15_21_0  (
            .in0(_gnd_net_),
            .in1(N__40804),
            .in2(N__40873),
            .in3(N__36764),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_15_21_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__47564),
            .ce(N__43567),
            .sr(N__46883));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_15_21_1  (
            .in0(_gnd_net_),
            .in1(N__41395),
            .in2(N__40838),
            .in3(N__36761),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__47564),
            .ce(N__43567),
            .sr(N__46883));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_15_21_2  (
            .in0(_gnd_net_),
            .in1(N__40805),
            .in2(N__41375),
            .in3(N__36758),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__47564),
            .ce(N__43567),
            .sr(N__46883));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_15_21_3  (
            .in0(_gnd_net_),
            .in1(N__41396),
            .in2(N__41216),
            .in3(N__36755),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__47564),
            .ce(N__43567),
            .sr(N__46883));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_15_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36752),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.T12_LC_15_23_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.T12_LC_15_23_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T12_LC_15_23_3 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \phase_controller_inst1.T12_LC_15_23_3  (
            .in0(N__36739),
            .in1(N__36579),
            .in2(_gnd_net_),
            .in3(N__36650),
            .lcout(T12_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47561),
            .ce(),
            .sr(N__46893));
    defparam \phase_controller_inst1.T45_LC_15_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.T45_LC_15_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T45_LC_15_24_4 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \phase_controller_inst1.T45_LC_15_24_4  (
            .in0(N__36710),
            .in1(N__38056),
            .in2(_gnd_net_),
            .in3(N__36721),
            .lcout(T45_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47559),
            .ce(),
            .sr(N__46898));
    defparam \phase_controller_inst1.T01_LC_15_24_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.T01_LC_15_24_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T01_LC_15_24_5 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \phase_controller_inst1.T01_LC_15_24_5  (
            .in0(N__36598),
            .in1(N__36709),
            .in2(_gnd_net_),
            .in3(N__36649),
            .lcout(T01_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47559),
            .ce(),
            .sr(N__46898));
    defparam \phase_controller_inst1.T23_LC_15_24_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.T23_LC_15_24_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.T23_LC_15_24_7 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \phase_controller_inst1.T23_LC_15_24_7  (
            .in0(N__36535),
            .in1(_gnd_net_),
            .in2(N__38060),
            .in3(N__36586),
            .lcout(T23_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47559),
            .ce(),
            .sr(N__46898));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_5_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_5_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_16_5_0  (
            .in0(N__38266),
            .in1(N__36889),
            .in2(_gnd_net_),
            .in3(N__48022),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_16_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_16_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_16_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_16_5_4  (
            .in0(N__38267),
            .in1(N__36888),
            .in2(_gnd_net_),
            .in3(N__48023),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47696),
            .ce(N__47209),
            .sr(N__46783));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_16_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_16_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_16_5_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_16_5_6  (
            .in0(N__38309),
            .in1(N__38097),
            .in2(_gnd_net_),
            .in3(N__48024),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47696),
            .ce(N__47209),
            .sr(N__46783));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_16_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_16_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_16_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_16_6_0  (
            .in0(N__48006),
            .in1(N__38118),
            .in2(_gnd_net_),
            .in3(N__38161),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47691),
            .ce(N__45955),
            .sr(N__46786));
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_16_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_16_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_16_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_21_LC_16_6_1  (
            .in0(N__41111),
            .in1(N__38414),
            .in2(_gnd_net_),
            .in3(N__48009),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47691),
            .ce(N__45955),
            .sr(N__46786));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_16_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_16_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_16_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_16_6_4  (
            .in0(N__48007),
            .in1(N__38301),
            .in2(_gnd_net_),
            .in3(N__38098),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47691),
            .ce(N__45955),
            .sr(N__46786));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_16_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_16_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_16_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_16_6_5  (
            .in0(N__41765),
            .in1(N__41738),
            .in2(_gnd_net_),
            .in3(N__48008),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47691),
            .ce(N__45955),
            .sr(N__46786));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_7_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_7_0  (
            .in0(N__36835),
            .in1(N__36785),
            .in2(N__36814),
            .in3(N__37016),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_16_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_16_7_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_16_7_1  (
            .in0(N__37015),
            .in1(N__36836),
            .in2(N__36815),
            .in3(N__36784),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_16_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_16_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_16_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_20_LC_16_7_2  (
            .in0(N__47995),
            .in1(N__38866),
            .in2(_gnd_net_),
            .in3(N__38911),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47680),
            .ce(N__45956),
            .sr(N__46789));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_16_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_16_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_16_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_16_7_4  (
            .in0(N__47996),
            .in1(N__38520),
            .in2(_gnd_net_),
            .in3(N__38498),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47680),
            .ce(N__45956),
            .sr(N__46789));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_16_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_16_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_16_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_16_7_6  (
            .in0(N__47997),
            .in1(N__41834),
            .in2(_gnd_net_),
            .in3(N__41809),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47680),
            .ce(N__45956),
            .sr(N__46789));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_16_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_16_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_16_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_16_7_7  (
            .in0(N__37040),
            .in1(N__37082),
            .in2(_gnd_net_),
            .in3(N__47998),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47680),
            .ce(N__45956),
            .sr(N__46789));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_16_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_16_8_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_16_8_0  (
            .in0(N__36976),
            .in1(N__36952),
            .in2(N__36917),
            .in3(N__36926),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_16_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_16_8_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_16_8_1  (
            .in0(N__36925),
            .in1(N__36977),
            .in2(N__36956),
            .in3(N__36913),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_16_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_16_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_16_8_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_22_LC_16_8_2  (
            .in0(N__48010),
            .in1(N__38558),
            .in2(_gnd_net_),
            .in3(N__41149),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47672),
            .ce(N__45957),
            .sr(N__46794));
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_16_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_16_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_16_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_23_LC_16_8_3  (
            .in0(N__48004),
            .in1(N__41692),
            .in2(_gnd_net_),
            .in3(N__41674),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47672),
            .ce(N__45957),
            .sr(N__46794));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_16_8_4  (
            .in0(N__37064),
            .in1(N__37097),
            .in2(_gnd_net_),
            .in3(N__48005),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47672),
            .ce(N__45957),
            .sr(N__46794));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_16_8_5  (
            .in0(N__48003),
            .in1(N__38698),
            .in2(_gnd_net_),
            .in3(N__38735),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47672),
            .ce(N__45957),
            .sr(N__46794));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_9_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_16_9_0  (
            .in0(N__37059),
            .in1(_gnd_net_),
            .in2(N__48179),
            .in3(N__37096),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_16_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_16_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_16_9_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__37060),
            .in2(N__37085),
            .in3(N__48096),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47659),
            .ce(N__47203),
            .sr(N__46800));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_16_9_2  (
            .in0(N__48091),
            .in1(N__37032),
            .in2(_gnd_net_),
            .in3(N__37078),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(elapsed_time_ns_1_RNIT6OBB_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_16_9_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_16_9_3  (
            .in0(N__37033),
            .in1(_gnd_net_),
            .in2(N__37067),
            .in3(N__48095),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47659),
            .ce(N__47203),
            .sr(N__46800));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_16_9_4  (
            .in0(N__37058),
            .in1(N__37031),
            .in2(N__38736),
            .in3(N__41791),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_16_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_16_9_7  (
            .in0(N__38738),
            .in1(N__38697),
            .in2(_gnd_net_),
            .in3(N__48097),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47659),
            .ce(N__47203),
            .sr(N__46800));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_10_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_16_10_0  (
            .in0(N__39053),
            .in1(N__38395),
            .in2(N__39077),
            .in3(N__37322),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_16_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_16_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_20_LC_16_10_2  (
            .in0(N__48099),
            .in1(N__38867),
            .in2(_gnd_net_),
            .in3(N__38903),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47649),
            .ce(N__47171),
            .sr(N__46808));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_10_3 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_16_10_3  (
            .in0(N__37321),
            .in1(N__39052),
            .in2(N__38399),
            .in3(N__39076),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_16_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_16_10_4  (
            .in0(N__48098),
            .in1(N__37313),
            .in2(_gnd_net_),
            .in3(N__37289),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47649),
            .ce(N__47171),
            .sr(N__46808));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_16_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_16_10_5  (
            .in0(N__38228),
            .in1(N__38192),
            .in2(_gnd_net_),
            .in3(N__48100),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47649),
            .ce(N__47171),
            .sr(N__46808));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_16_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_16_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_16_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_16_10_7  (
            .in0(N__37247),
            .in1(N__37220),
            .in2(_gnd_net_),
            .in3(N__48101),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47649),
            .ce(N__47171),
            .sr(N__46808));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_16_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_16_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__37184),
            .in2(N__37193),
            .in3(N__38670),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_16_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_16_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__37178),
            .in2(N__37172),
            .in3(N__38647),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_16_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_16_11_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_16_11_2  (
            .in0(N__38632),
            .in1(N__37163),
            .in2(N__37151),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_16_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_16_11_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_16_11_3  (
            .in0(N__38617),
            .in1(N__37133),
            .in2(N__37142),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_16_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_16_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__37127),
            .in2(N__37115),
            .in3(N__39031),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_16_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_16_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_16_11_5  (
            .in0(N__39016),
            .in1(N__37433),
            .in2(N__37424),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_16_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_16_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_16_11_6  (
            .in0(N__39001),
            .in1(N__38534),
            .in2(N__37415),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_16_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_16_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(N__37406),
            .in2(N__38471),
            .in3(N__38986),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_16_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_16_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__37400),
            .in2(N__41780),
            .in3(N__38971),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_16_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_16_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__37382),
            .in2(N__37394),
            .in3(N__38956),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_16_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_16_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__37376),
            .in2(N__37367),
            .in3(N__38941),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_16_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_16_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__37358),
            .in2(N__37349),
            .in3(N__38926),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_16_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_16_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_16_12_4  (
            .in0(N__39133),
            .in1(N__37328),
            .in2(N__37340),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_16_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_16_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_16_12_5  (
            .in0(N__39118),
            .in1(N__41471),
            .in2(N__37478),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_16_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_16_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(N__42488),
            .in2(N__37466),
            .in3(N__39103),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_16_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_16_12_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(N__41540),
            .in2(N__41618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_16_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_16_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__41996),
            .in2(N__41951),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_16_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_16_13_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__37457),
            .in2(N__37448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_16_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_16_13_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__38588),
            .in2(N__38573),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_16_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_16_13_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__46379),
            .in2(N__46460),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_16_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_16_13_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__45566),
            .in2(N__46295),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_16_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_16_13_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__45647),
            .in2(N__45578),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_LUT4_0_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__42110),
            .in2(N__37526),
            .in3(N__37511),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_28_THRU_CO ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37508),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_16_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_16_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__45079),
            .in2(N__37505),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_16_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_16_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__37947),
            .in2(N__37487),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_16_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_16_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__39293),
            .in2(N__37994),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_16_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_16_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(N__37951),
            .in2(N__39248),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_16_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_16_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__39380),
            .in2(N__37995),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_16_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_16_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(N__37955),
            .in2(N__39788),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_16_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_16_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__39287),
            .in2(N__37996),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_16_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_16_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(N__37959),
            .in2(N__39335),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_16_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_16_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__37943),
            .in2(N__39416),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_16_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_16_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__39458),
            .in2(N__37993),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_16_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_16_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__37931),
            .in2(N__39629),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_16_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_16_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__39578),
            .in2(N__37990),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_16_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_16_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__37935),
            .in2(N__39674),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_16_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_16_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__39716),
            .in2(N__37991),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_16_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_16_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__37939),
            .in2(N__39779),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_16_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_16_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__39536),
            .in2(N__37992),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_16_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_16_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__37761),
            .in2(N__40082),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_16_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_16_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__39977),
            .in2(N__37843),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_16_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_16_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__37765),
            .in2(N__39887),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_16_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_16_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__37532),
            .in2(N__37844),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_16_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_16_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__37769),
            .in2(N__39842),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_16_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_16_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(N__39932),
            .in2(N__37845),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_16_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_16_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(N__37773),
            .in2(N__39986),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_16_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_16_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(N__39938),
            .in2(N__37846),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_16_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_16_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__40310),
            .in2(N__37997),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_16_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_16_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(N__37963),
            .in2(N__40031),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_16_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_16_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(N__40160),
            .in2(N__37998),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_16_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_16_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(N__37967),
            .in2(N__40277),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_16_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_16_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__40268),
            .in2(N__37999),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_16_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_16_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(N__37971),
            .in2(N__39833),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_16_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_16_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(N__43694),
            .in2(N__38000),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_17_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(N__44390),
            .in2(_gnd_net_),
            .in3(N__37637),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_18_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__39266),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39391),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39804),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__39306),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39687),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40095),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39552),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39999),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_16_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_16_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNI7NN7_LC_16_19_4  (
            .in0(N__38081),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38055),
            .lcout(\phase_controller_inst1.time_passed_RNI7NN7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_19_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42444),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39727),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_16_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_16_20_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39951),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_16_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40288),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39900),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_16_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39860),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_16_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40328),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40178),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_21_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40248),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_17_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_17_5_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_17_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_17_5_1  (
            .in0(N__38184),
            .in1(N__38227),
            .in2(_gnd_net_),
            .in3(N__48019),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_17_5_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_17_5_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_17_5_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_17_5_6  (
            .in0(N__48020),
            .in1(N__38119),
            .in2(_gnd_net_),
            .in3(N__38165),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_17_5_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_17_5_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_17_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_17_5_7  (
            .in0(N__38099),
            .in1(N__38308),
            .in2(_gnd_net_),
            .in3(N__48021),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_17_6_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_17_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_17_6_3  (
            .in0(N__41906),
            .in1(N__42596),
            .in2(N__41741),
            .in3(N__38912),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_17_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_17_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_17_6_5  (
            .in0(N__41113),
            .in1(N__38413),
            .in2(_gnd_net_),
            .in3(N__47986),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(elapsed_time_ns_1_RNIV9PBB_0_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_17_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_17_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_17_6_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_21_LC_17_6_6  (
            .in0(N__47987),
            .in1(_gnd_net_),
            .in2(N__38402),
            .in3(N__41114),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47697),
            .ce(N__47229),
            .sr(N__46784));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_17_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_17_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_17_7_0  (
            .in0(N__41069),
            .in1(N__41024),
            .in2(N__38381),
            .in3(N__38423),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_17_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_17_7_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_17_7_1  (
            .in0(N__45704),
            .in1(N__48284),
            .in2(_gnd_net_),
            .in3(N__38369),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_2 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_17_7_2  (
            .in0(N__38357),
            .in1(N__38594),
            .in2(N__38321),
            .in3(N__38318),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_17_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_17_7_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(N__38500),
            .in2(N__38312),
            .in3(N__38521),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_17_7_4  (
            .in0(N__38499),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38795),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_17_7_5  (
            .in0(N__38300),
            .in1(N__38264),
            .in2(N__38231),
            .in3(N__38603),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_17_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_17_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_17_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_17_7_7  (
            .in0(N__41693),
            .in1(N__41673),
            .in2(_gnd_net_),
            .in3(N__47988),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_8_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_17_8_0  (
            .in0(N__39235),
            .in1(N__41630),
            .in2(N__39212),
            .in3(N__38543),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_17_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_17_8_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_17_8_1  (
            .in0(N__38542),
            .in1(N__39208),
            .in2(N__39239),
            .in3(N__41629),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_17_8_4  (
            .in0(N__41147),
            .in1(N__38557),
            .in2(_gnd_net_),
            .in3(N__47982),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_17_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_17_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_17_8_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_22_LC_17_8_5  (
            .in0(N__47983),
            .in1(_gnd_net_),
            .in2(N__38546),
            .in3(N__41148),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47681),
            .ce(N__47220),
            .sr(N__46790));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_17_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_17_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_17_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_17_8_6  (
            .in0(N__38754),
            .in1(N__38797),
            .in2(_gnd_net_),
            .in3(N__47985),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47681),
            .ce(N__47220),
            .sr(N__46790));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_17_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_17_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_17_8_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_17_8_7  (
            .in0(N__47984),
            .in1(_gnd_net_),
            .in2(N__38522),
            .in3(N__38501),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47681),
            .ce(N__47220),
            .sr(N__46790));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_17_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_17_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_17_9_0  (
            .in0(N__42546),
            .in1(N__41501),
            .in2(N__38459),
            .in3(N__41447),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_17_9_1  (
            .in0(N__42510),
            .in1(N__42547),
            .in2(_gnd_net_),
            .in3(N__48087),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_17_9_2  (
            .in0(N__48089),
            .in1(N__38865),
            .in2(_gnd_net_),
            .in3(N__38910),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_17_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_17_9_3 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_RNI42MA1_30_LC_17_9_3  (
            .in0(N__39165),
            .in1(N__38846),
            .in2(N__39527),
            .in3(N__38825),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_df30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_17_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_17_9_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_17_9_4  (
            .in0(N__48088),
            .in1(N__38758),
            .in2(_gnd_net_),
            .in3(N__38796),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_17_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_17_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_17_9_5  (
            .in0(N__38699),
            .in1(N__38737),
            .in2(_gnd_net_),
            .in3(N__48090),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__42002),
            .in2(N__38681),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_17_10_1  (
            .in0(N__47113),
            .in1(N__38648),
            .in2(_gnd_net_),
            .in3(N__38636),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__47660),
            .ce(),
            .sr(N__46801));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_10_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_17_10_2  (
            .in0(N__47117),
            .in1(N__38633),
            .in2(N__42158),
            .in3(N__38621),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__47660),
            .ce(),
            .sr(N__46801));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_17_10_3  (
            .in0(N__47114),
            .in1(N__38618),
            .in2(_gnd_net_),
            .in3(N__38606),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__47660),
            .ce(),
            .sr(N__46801));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_17_10_4  (
            .in0(N__47118),
            .in1(N__39032),
            .in2(_gnd_net_),
            .in3(N__39020),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__47660),
            .ce(),
            .sr(N__46801));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_17_10_5  (
            .in0(N__47115),
            .in1(N__39017),
            .in2(_gnd_net_),
            .in3(N__39005),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__47660),
            .ce(),
            .sr(N__46801));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_17_10_6  (
            .in0(N__47119),
            .in1(N__39002),
            .in2(_gnd_net_),
            .in3(N__38990),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__47660),
            .ce(),
            .sr(N__46801));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_17_10_7  (
            .in0(N__47116),
            .in1(N__38987),
            .in2(_gnd_net_),
            .in3(N__38975),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__47660),
            .ce(),
            .sr(N__46801));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_17_11_0  (
            .in0(N__47157),
            .in1(N__38972),
            .in2(_gnd_net_),
            .in3(N__38960),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__47650),
            .ce(),
            .sr(N__46809));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_17_11_1  (
            .in0(N__47150),
            .in1(N__38957),
            .in2(_gnd_net_),
            .in3(N__38945),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__47650),
            .ce(),
            .sr(N__46809));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_17_11_2  (
            .in0(N__47154),
            .in1(N__38942),
            .in2(_gnd_net_),
            .in3(N__38930),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__47650),
            .ce(),
            .sr(N__46809));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_17_11_3  (
            .in0(N__47151),
            .in1(N__38927),
            .in2(_gnd_net_),
            .in3(N__38915),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__47650),
            .ce(),
            .sr(N__46809));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_17_11_4  (
            .in0(N__47155),
            .in1(N__39134),
            .in2(_gnd_net_),
            .in3(N__39122),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__47650),
            .ce(),
            .sr(N__46809));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_17_11_5  (
            .in0(N__47152),
            .in1(N__39119),
            .in2(_gnd_net_),
            .in3(N__39107),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__47650),
            .ce(),
            .sr(N__46809));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_17_11_6  (
            .in0(N__47156),
            .in1(N__39104),
            .in2(_gnd_net_),
            .in3(N__39092),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__47650),
            .ce(),
            .sr(N__46809));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_17_11_7  (
            .in0(N__47153),
            .in1(N__41587),
            .in2(_gnd_net_),
            .in3(N__39089),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__47650),
            .ce(),
            .sr(N__46809));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_17_12_0  (
            .in0(N__47158),
            .in1(N__41568),
            .in2(_gnd_net_),
            .in3(N__39086),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__47637),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_17_12_1  (
            .in0(N__47162),
            .in1(N__41968),
            .in2(_gnd_net_),
            .in3(N__39083),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__47637),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_17_12_2  (
            .in0(N__47159),
            .in1(N__41984),
            .in2(_gnd_net_),
            .in3(N__39080),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__47637),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_17_12_3  (
            .in0(N__47163),
            .in1(N__39072),
            .in2(_gnd_net_),
            .in3(N__39056),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__47637),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_17_12_4  (
            .in0(N__47160),
            .in1(N__39051),
            .in2(_gnd_net_),
            .in3(N__39035),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__47637),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_17_12_5  (
            .in0(N__47164),
            .in1(N__39234),
            .in2(_gnd_net_),
            .in3(N__39215),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__47637),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_17_12_6  (
            .in0(N__47161),
            .in1(N__39207),
            .in2(_gnd_net_),
            .in3(N__39191),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__47637),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_17_12_7  (
            .in0(N__47165),
            .in1(N__46402),
            .in2(_gnd_net_),
            .in3(N__39188),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__47637),
            .ce(),
            .sr(N__46818));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_17_13_0  (
            .in0(N__47067),
            .in1(N__46434),
            .in2(_gnd_net_),
            .in3(N__39185),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__47627),
            .ce(),
            .sr(N__46828));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_17_13_1  (
            .in0(N__47188),
            .in1(N__46365),
            .in2(_gnd_net_),
            .in3(N__39182),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__47627),
            .ce(),
            .sr(N__46828));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_17_13_2  (
            .in0(N__47068),
            .in1(N__46329),
            .in2(_gnd_net_),
            .in3(N__39179),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__47627),
            .ce(),
            .sr(N__46828));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_17_13_3  (
            .in0(N__47189),
            .in1(N__45615),
            .in2(_gnd_net_),
            .in3(N__39176),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__47627),
            .ce(),
            .sr(N__46828));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_17_13_4  (
            .in0(N__47069),
            .in1(N__45594),
            .in2(_gnd_net_),
            .in3(N__39173),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__47627),
            .ce(),
            .sr(N__46828));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_17_13_5  (
            .in0(N__47190),
            .in1(N__39159),
            .in2(_gnd_net_),
            .in3(N__39137),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__47627),
            .ce(),
            .sr(N__46828));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_17_13_6  (
            .in0(N__47070),
            .in1(N__39516),
            .in2(_gnd_net_),
            .in3(N__39530),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47627),
            .ce(),
            .sr(N__46828));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_14_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_17_14_0  (
            .in0(N__42313),
            .in1(N__39494),
            .in2(_gnd_net_),
            .in3(N__42702),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_14_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_17_14_1  (
            .in0(N__42317),
            .in1(N__39452),
            .in2(_gnd_net_),
            .in3(N__42747),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_17_14_2  (
            .in0(N__42312),
            .in1(N__39405),
            .in2(_gnd_net_),
            .in3(N__42876),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_17_14_3  (
            .in0(N__42316),
            .in1(N__39369),
            .in2(_gnd_net_),
            .in3(N__42792),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_14_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_17_14_4  (
            .in0(N__42310),
            .in1(N__39321),
            .in2(_gnd_net_),
            .in3(N__42217),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_17_14_5  (
            .in0(N__42315),
            .in1(N__43685),
            .in2(_gnd_net_),
            .in3(N__43644),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_17_14_6  (
            .in0(N__42311),
            .in1(N__39280),
            .in2(_gnd_net_),
            .in3(N__42177),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_14_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_17_14_7  (
            .in0(N__42314),
            .in1(N__39822),
            .in2(_gnd_net_),
            .in3(N__42838),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_15_0  (
            .in0(N__44062),
            .in1(N__42362),
            .in2(_gnd_net_),
            .in3(N__43101),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_17_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_17_15_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNO_LC_17_15_1  (
            .in0(N__43680),
            .in1(N__44418),
            .in2(N__45038),
            .in3(N__43645),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_15_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_15_2  (
            .in0(N__39750),
            .in1(N__42361),
            .in2(_gnd_net_),
            .in3(N__43140),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_15_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_17_15_3  (
            .in0(N__42360),
            .in1(N__39702),
            .in2(_gnd_net_),
            .in3(N__43177),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43679),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_17_15_5  (
            .in0(N__42358),
            .in1(N__39660),
            .in2(_gnd_net_),
            .in3(N__42660),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_15_6  (
            .in0(N__39615),
            .in1(N__42359),
            .in2(_gnd_net_),
            .in3(N__42621),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_17_15_7  (
            .in0(N__42363),
            .in1(N__39572),
            .in2(_gnd_net_),
            .in3(N__43062),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_17_16_0  (
            .in0(N__40113),
            .in1(N__42364),
            .in2(_gnd_net_),
            .in3(N__43017),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_17_16_1  (
            .in0(N__44426),
            .in1(N__40073),
            .in2(_gnd_net_),
            .in3(N__43290),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_16_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_17_16_2  (
            .in0(N__40017),
            .in1(N__42369),
            .in2(_gnd_net_),
            .in3(N__43423),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_17_16_3  (
            .in0(N__42365),
            .in1(_gnd_net_),
            .in2(N__42994),
            .in3(N__43959),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_4 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_17_16_4  (
            .in0(N__43392),
            .in1(N__39969),
            .in2(_gnd_net_),
            .in3(N__42370),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_16_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_17_16_5  (
            .in0(N__42368),
            .in1(N__42462),
            .in2(_gnd_net_),
            .in3(N__43473),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_16_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_17_16_6  (
            .in0(N__39918),
            .in1(N__42366),
            .in2(_gnd_net_),
            .in3(N__42948),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_17_16_7  (
            .in0(N__42367),
            .in1(N__39877),
            .in2(_gnd_net_),
            .in3(N__43506),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_17_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_17_17_0  (
            .in0(N__44007),
            .in1(N__44424),
            .in2(_gnd_net_),
            .in3(N__43716),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_17_17_1  (
            .in0(N__42382),
            .in1(N__40347),
            .in2(_gnd_net_),
            .in3(N__43341),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_17_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_17_17_2  (
            .in0(N__44427),
            .in1(N__40302),
            .in2(_gnd_net_),
            .in3(N__43210),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_17_17_3  (
            .in0(N__44423),
            .in1(N__40261),
            .in2(_gnd_net_),
            .in3(N__43743),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_4 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_17_17_4  (
            .in0(N__40262),
            .in1(N__44425),
            .in2(N__43750),
            .in3(N__44961),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_17_5  (
            .in0(N__44421),
            .in1(N__42466),
            .in2(N__45039),
            .in3(N__43474),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_17_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNO_LC_17_17_6  (
            .in0(N__44965),
            .in1(N__44420),
            .in2(N__43966),
            .in3(N__42993),
            .lcout(\current_shift_inst.un38_control_input_cry_17_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_17_17_7  (
            .in0(N__44422),
            .in1(N__40193),
            .in2(_gnd_net_),
            .in3(N__43248),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_17_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_17_18_0  (
            .in0(N__41325),
            .in1(N__40146),
            .in2(_gnd_net_),
            .in3(N__40127),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__47582),
            .ce(N__41197),
            .sr(N__46858));
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_17_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_17_18_1  (
            .in0(N__41351),
            .in1(N__43593),
            .in2(_gnd_net_),
            .in3(N__40124),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__47582),
            .ce(N__41197),
            .sr(N__46858));
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_17_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_17_18_2  (
            .in0(N__41326),
            .in1(N__40566),
            .in2(_gnd_net_),
            .in3(N__40550),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__47582),
            .ce(N__41197),
            .sr(N__46858));
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_17_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_17_18_3  (
            .in0(N__41352),
            .in1(N__40536),
            .in2(_gnd_net_),
            .in3(N__40520),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__47582),
            .ce(N__41197),
            .sr(N__46858));
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_17_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_17_18_4  (
            .in0(N__41327),
            .in1(N__40509),
            .in2(_gnd_net_),
            .in3(N__40493),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__47582),
            .ce(N__41197),
            .sr(N__46858));
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_17_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_17_18_5  (
            .in0(N__41353),
            .in1(N__40482),
            .in2(_gnd_net_),
            .in3(N__40466),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__47582),
            .ce(N__41197),
            .sr(N__46858));
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_17_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_17_18_6  (
            .in0(N__41328),
            .in1(N__40461),
            .in2(_gnd_net_),
            .in3(N__40445),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__47582),
            .ce(N__41197),
            .sr(N__46858));
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_17_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_17_18_7  (
            .in0(N__41354),
            .in1(N__40440),
            .in2(_gnd_net_),
            .in3(N__40424),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__47582),
            .ce(N__41197),
            .sr(N__46858));
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_17_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_17_19_0  (
            .in0(N__41344),
            .in1(N__40413),
            .in2(_gnd_net_),
            .in3(N__40391),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__47578),
            .ce(N__41198),
            .sr(N__46863));
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_17_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_17_19_1  (
            .in0(N__41340),
            .in1(N__40374),
            .in2(_gnd_net_),
            .in3(N__40355),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__47578),
            .ce(N__41198),
            .sr(N__46863));
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_17_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_17_19_2  (
            .in0(N__41341),
            .in1(N__40782),
            .in2(_gnd_net_),
            .in3(N__40766),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__47578),
            .ce(N__41198),
            .sr(N__46863));
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_17_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_17_19_3  (
            .in0(N__41337),
            .in1(N__40761),
            .in2(_gnd_net_),
            .in3(N__40745),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__47578),
            .ce(N__41198),
            .sr(N__46863));
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_17_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_17_19_4  (
            .in0(N__41342),
            .in1(N__40737),
            .in2(_gnd_net_),
            .in3(N__40718),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__47578),
            .ce(N__41198),
            .sr(N__46863));
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_17_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_17_19_5  (
            .in0(N__41338),
            .in1(N__40710),
            .in2(_gnd_net_),
            .in3(N__40691),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__47578),
            .ce(N__41198),
            .sr(N__46863));
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_17_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_17_19_6  (
            .in0(N__41343),
            .in1(N__40680),
            .in2(_gnd_net_),
            .in3(N__40664),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__47578),
            .ce(N__41198),
            .sr(N__46863));
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_17_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_17_19_7  (
            .in0(N__41339),
            .in1(N__40653),
            .in2(_gnd_net_),
            .in3(N__40637),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__47578),
            .ce(N__41198),
            .sr(N__46863));
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_17_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_17_20_0  (
            .in0(N__41347),
            .in1(N__40626),
            .in2(_gnd_net_),
            .in3(N__40604),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__47573),
            .ce(N__41193),
            .sr(N__46868));
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_17_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_17_20_1  (
            .in0(N__41333),
            .in1(N__40587),
            .in2(_gnd_net_),
            .in3(N__40571),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__47573),
            .ce(N__41193),
            .sr(N__46868));
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_17_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_17_20_2  (
            .in0(N__41348),
            .in1(N__41016),
            .in2(_gnd_net_),
            .in3(N__41000),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__47573),
            .ce(N__41193),
            .sr(N__46868));
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_17_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_17_20_3  (
            .in0(N__41334),
            .in1(N__40992),
            .in2(_gnd_net_),
            .in3(N__40973),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__47573),
            .ce(N__41193),
            .sr(N__46868));
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_17_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_17_20_4  (
            .in0(N__41349),
            .in1(N__40962),
            .in2(_gnd_net_),
            .in3(N__40946),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__47573),
            .ce(N__41193),
            .sr(N__46868));
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_17_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_17_20_5  (
            .in0(N__41335),
            .in1(N__40941),
            .in2(_gnd_net_),
            .in3(N__40925),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__47573),
            .ce(N__41193),
            .sr(N__46868));
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_17_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_17_20_6  (
            .in0(N__41350),
            .in1(N__40920),
            .in2(_gnd_net_),
            .in3(N__40904),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__47573),
            .ce(N__41193),
            .sr(N__46868));
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_17_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_17_20_7  (
            .in0(N__41336),
            .in1(N__40893),
            .in2(_gnd_net_),
            .in3(N__40877),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__47573),
            .ce(N__41193),
            .sr(N__46868));
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_17_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_17_21_0  (
            .in0(N__41329),
            .in1(N__40863),
            .in2(_gnd_net_),
            .in3(N__40841),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__47568),
            .ce(N__41186),
            .sr(N__46872));
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_17_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_17_21_1  (
            .in0(N__41345),
            .in1(N__40830),
            .in2(_gnd_net_),
            .in3(N__40808),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__47568),
            .ce(N__41186),
            .sr(N__46872));
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_17_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_17_21_2  (
            .in0(N__41330),
            .in1(N__40803),
            .in2(_gnd_net_),
            .in3(N__40787),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__47568),
            .ce(N__41186),
            .sr(N__46872));
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_17_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_17_21_3  (
            .in0(N__41346),
            .in1(N__41394),
            .in2(_gnd_net_),
            .in3(N__41378),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__47568),
            .ce(N__41186),
            .sr(N__46872));
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_17_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_17_21_4  (
            .in0(N__41331),
            .in1(N__41371),
            .in2(_gnd_net_),
            .in3(N__41357),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__47568),
            .ce(N__41186),
            .sr(N__46872));
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_17_21_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_17_21_5  (
            .in0(N__41212),
            .in1(N__41332),
            .in2(_gnd_net_),
            .in3(N__41219),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47568),
            .ce(N__41186),
            .sr(N__46872));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_18_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_18_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_18_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_18_6_4  (
            .in0(N__41672),
            .in1(N__41150),
            .in2(N__45840),
            .in3(N__41112),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_18_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_18_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_18_7_1  (
            .in0(N__41764),
            .in1(N__41739),
            .in2(_gnd_net_),
            .in3(N__47980),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_18_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_18_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_18_7_2  (
            .in0(N__45926),
            .in1(N__45757),
            .in2(N__47777),
            .in3(N__41062),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_18_7_7  (
            .in0(N__41833),
            .in1(N__41808),
            .in2(_gnd_net_),
            .in3(N__47981),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_18_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_18_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_18_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_18_8_0  (
            .in0(N__41459),
            .in1(N__41416),
            .in2(_gnd_net_),
            .in3(N__48001),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47692),
            .ce(N__47204),
            .sr(N__46787));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_18_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_18_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_18_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_18_8_5  (
            .in0(N__48000),
            .in1(N__41829),
            .in2(_gnd_net_),
            .in3(N__41813),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47692),
            .ce(N__47204),
            .sr(N__46787));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_18_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_18_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_18_8_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_18_8_6  (
            .in0(N__41754),
            .in1(_gnd_net_),
            .in2(N__41740),
            .in3(N__48002),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47692),
            .ce(N__47204),
            .sr(N__46787));
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_18_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_18_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_18_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_23_LC_18_8_7  (
            .in0(N__47999),
            .in1(N__41691),
            .in2(_gnd_net_),
            .in3(N__41675),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47692),
            .ce(N__47204),
            .sr(N__46787));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_18_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_18_9_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_18_9_0  (
            .in0(N__41593),
            .in1(N__41603),
            .in2(N__41552),
            .in3(N__41572),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_18_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_18_9_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_18_9_1  (
            .in0(N__41602),
            .in1(N__41594),
            .in2(N__41573),
            .in3(N__41551),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_18_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_18_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_18_9_6  (
            .in0(N__41528),
            .in1(N__41502),
            .in2(_gnd_net_),
            .in3(N__48051),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47682),
            .ce(N__47202),
            .sr(N__46791));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_18_10_0  (
            .in0(N__41415),
            .in1(N__41455),
            .in2(_gnd_net_),
            .in3(N__48026),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_10_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_18_10_1  (
            .in0(N__48025),
            .in1(N__41925),
            .in2(_gnd_net_),
            .in3(N__41905),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_18_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_18_10_4 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_18_10_4  (
            .in0(N__45497),
            .in1(N__42121),
            .in2(_gnd_net_),
            .in3(N__45556),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(\phase_controller_inst1.stoper_tr.un2_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_18_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_18_10_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4_28_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42161),
            .in3(N__42058),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIO3KK4Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_LC_18_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_18_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_18_11_3 .LUT_INIT=16'b1101010111001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_18_11_3  (
            .in0(N__45499),
            .in1(N__42122),
            .in2(N__42149),
            .in3(N__42021),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47661),
            .ce(),
            .sr(N__46802));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_18_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_18_11_4 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNIIMJC3_28_LC_18_11_4  (
            .in0(N__42109),
            .in1(N__45498),
            .in2(N__42086),
            .in3(N__42074),
            .lcout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i ),
            .ltout(\phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_11_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42047),
            .in3(N__42020),
            .lcout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_12_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_18_12_0  (
            .in0(N__41982),
            .in1(N__41964),
            .in2(N__41867),
            .in3(N__42560),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_18_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_18_12_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_18_12_1  (
            .in0(N__42559),
            .in1(N__41983),
            .in2(N__41969),
            .in3(N__41863),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_18_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_18_12_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_18_12_3  (
            .in0(N__48131),
            .in1(_gnd_net_),
            .in2(N__41935),
            .in3(N__41900),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47651),
            .ce(N__47172),
            .sr(N__46810));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_12_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_18_12_4  (
            .in0(N__42597),
            .in1(N__41845),
            .in2(_gnd_net_),
            .in3(N__48129),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(elapsed_time_ns_1_RNI5FOBB_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_18_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_18_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_18_12_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_18_12_5  (
            .in0(N__48130),
            .in1(_gnd_net_),
            .in2(N__42602),
            .in3(N__42598),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47651),
            .ce(N__47172),
            .sr(N__46810));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_18_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_18_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_18_12_6  (
            .in0(N__42551),
            .in1(N__42517),
            .in2(_gnd_net_),
            .in3(N__48132),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47651),
            .ce(N__47172),
            .sr(N__46810));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_13_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_13_3  (
            .in0(N__44415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44954),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_13_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_18_13_4  (
            .in0(N__42467),
            .in1(N__44414),
            .in2(N__45037),
            .in3(N__43478),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42414),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47638),
            .ce(N__43574),
            .sr(N__46819));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_18_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_18_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__43544),
            .in2(N__42266),
            .in3(N__42265),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_18_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_18_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__42242),
            .in2(_gnd_net_),
            .in3(N__42206),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_18_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_18_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__42203),
            .in2(_gnd_net_),
            .in3(N__42164),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_18_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_18_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__42902),
            .in2(_gnd_net_),
            .in3(N__42863),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_18_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_18_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__42860),
            .in2(_gnd_net_),
            .in3(N__42827),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_18_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_18_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__42824),
            .in2(_gnd_net_),
            .in3(N__42818),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_18_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_18_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__42815),
            .in2(_gnd_net_),
            .in3(N__42776),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_18_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_18_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__42773),
            .in2(_gnd_net_),
            .in3(N__42734),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_18_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_18_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__42731),
            .in2(_gnd_net_),
            .in3(N__42689),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_18_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_18_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(N__42686),
            .in2(_gnd_net_),
            .in3(N__42647),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_18_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_18_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(N__42644),
            .in2(_gnd_net_),
            .in3(N__42605),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_18_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_18_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_18_15_3  (
            .in0(_gnd_net_),
            .in1(N__43196),
            .in2(_gnd_net_),
            .in3(N__43166),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_18_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_18_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__43163),
            .in2(_gnd_net_),
            .in3(N__43124),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_18_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_18_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(N__44024),
            .in2(_gnd_net_),
            .in3(N__43085),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_18_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_18_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__43082),
            .in2(_gnd_net_),
            .in3(N__43046),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_18_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_18_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__43043),
            .in2(_gnd_net_),
            .in3(N__43001),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_18_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_18_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__43916),
            .in2(_gnd_net_),
            .in3(N__42971),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_18_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_18_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__42968),
            .in2(_gnd_net_),
            .in3(N__42935),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_18_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_18_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__43871),
            .in2(_gnd_net_),
            .in3(N__42905),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_18_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_18_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__43532),
            .in2(_gnd_net_),
            .in3(N__43493),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_18_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_18_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(N__43490),
            .in2(_gnd_net_),
            .in3(N__43457),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_18_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_18_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__43454),
            .in2(_gnd_net_),
            .in3(N__43412),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_18_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_18_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__43409),
            .in2(_gnd_net_),
            .in3(N__43370),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_18_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_18_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(N__43367),
            .in2(_gnd_net_),
            .in3(N__43325),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_18_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_18_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__43322),
            .in2(_gnd_net_),
            .in3(N__43277),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_18_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_18_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__43274),
            .in2(_gnd_net_),
            .in3(N__43232),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_18_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_18_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__43229),
            .in2(_gnd_net_),
            .in3(N__43199),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_18_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_18_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__43766),
            .in2(_gnd_net_),
            .in3(N__43730),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_18_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_18_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__43976),
            .in2(_gnd_net_),
            .in3(N__43703),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_18_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_18_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43700),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(\current_shift_inst.un4_control_input1_31_THRU_CO_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_17_6 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43697),
            .in3(N__44397),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_18_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_18_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNO_LC_18_17_7  (
            .in0(N__44396),
            .in1(N__43684),
            .in2(N__45055),
            .in3(N__43649),
            .lcout(\current_shift_inst.un38_control_input_cry_6_s0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_18_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_18_18_0  (
            .in0(N__44393),
            .in1(N__45218),
            .in2(N__45167),
            .in3(N__45186),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43594),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47588),
            .ce(N__43573),
            .sr(N__46852));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45182),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_18_3 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_18_3  (
            .in0(N__45217),
            .in1(N__44392),
            .in2(N__45190),
            .in3(N__45166),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_18_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_18_18_6  (
            .in0(N__44394),
            .in1(N__45050),
            .in2(N__45092),
            .in3(N__45100),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_18_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_18_18_7  (
            .in0(N__45101),
            .in1(N__45088),
            .in2(N__45056),
            .in3(N__44395),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_19_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44046),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_18_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_18_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43997),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_19_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43949),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_18_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_18_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43890),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_18_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_18_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_18_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43862),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47566),
            .ce(),
            .sr(N__46877));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_9_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_20_9_0  (
            .in0(N__45418),
            .in1(N__45971),
            .in2(N__45449),
            .in3(N__45992),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_9_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_20_9_1  (
            .in0(N__45991),
            .in1(N__45448),
            .in2(N__45422),
            .in3(N__45970),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_20_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_20_9_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_20_9_4  (
            .in0(N__45310),
            .in1(N__45371),
            .in2(N__45347),
            .in3(N__45979),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_9_5 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_9_5  (
            .in0(N__45370),
            .in1(N__45311),
            .in2(N__45983),
            .in3(N__45346),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_20_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_20_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_20_9_7  (
            .in0(N__45705),
            .in1(N__45667),
            .in2(_gnd_net_),
            .in3(N__48152),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_20_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_20_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_20_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_26_LC_20_10_0  (
            .in0(N__45787),
            .in1(N__45770),
            .in2(_gnd_net_),
            .in3(N__48178),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47693),
            .ce(N__45958),
            .sr(N__46795));
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_20_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_20_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_20_10_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_29_LC_20_10_1  (
            .in0(N__48177),
            .in1(N__45884),
            .in2(_gnd_net_),
            .in3(N__45928),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47693),
            .ce(N__45958),
            .sr(N__46795));
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_20_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_20_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_20_10_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_28_LC_20_10_3  (
            .in0(N__48176),
            .in1(N__45713),
            .in2(_gnd_net_),
            .in3(N__45663),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47693),
            .ce(N__45958),
            .sr(N__46795));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_11_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_11_0  (
            .in0(N__45227),
            .in1(N__45287),
            .in2(N__45256),
            .in3(N__45278),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_20_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_20_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_20_11_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_20_11_1  (
            .in0(N__45286),
            .in1(N__45277),
            .in2(N__45257),
            .in3(N__45226),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_20_11_2  (
            .in0(N__47722),
            .in1(N__48151),
            .in2(_gnd_net_),
            .in3(N__47775),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_20_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_20_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_20_12_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_28_LC_20_12_0  (
            .in0(N__45712),
            .in1(N__45668),
            .in2(_gnd_net_),
            .in3(N__48199),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47674),
            .ce(N__47237),
            .sr(N__46811));
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_29_LC_20_12_3  (
            .in0(N__48198),
            .in1(N__45883),
            .in2(_gnd_net_),
            .in3(N__45929),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47674),
            .ce(N__47237),
            .sr(N__46811));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_20_13_0  (
            .in0(_gnd_net_),
            .in1(N__45488),
            .in2(_gnd_net_),
            .in3(N__45557),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_20_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_20_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_20_13_4 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_20_13_4  (
            .in0(N__45628),
            .in1(N__45619),
            .in2(N__45599),
            .in3(N__45637),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_13_5 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_20_13_5  (
            .in0(N__45638),
            .in1(N__45629),
            .in2(N__45620),
            .in3(N__45598),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_13_7 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_20_13_7  (
            .in0(N__46346),
            .in1(N__46330),
            .in2(N__46370),
            .in3(N__46307),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_20_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_20_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_20_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_20_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45555),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47640),
            .ce(),
            .sr(N__46834));
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_21_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_21_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_21_9_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_24_LC_21_9_3  (
            .in0(N__45863),
            .in1(_gnd_net_),
            .in2(N__48204),
            .in3(N__45842),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47700),
            .ce(N__45959),
            .sr(N__46796));
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_21_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_21_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_21_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_27_LC_21_9_4  (
            .in0(N__48286),
            .in1(N__48169),
            .in2(_gnd_net_),
            .in3(N__48222),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47700),
            .ce(N__45959),
            .sr(N__46796));
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_21_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_21_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_21_9_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_25_LC_21_9_7  (
            .in0(N__47723),
            .in1(_gnd_net_),
            .in2(N__48205),
            .in3(N__47776),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47700),
            .ce(N__45959),
            .sr(N__46796));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_21_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_21_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_21_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_21_10_0  (
            .in0(N__48285),
            .in1(N__48226),
            .in2(_gnd_net_),
            .in3(N__48153),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_21_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_21_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_21_10_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_21_10_1  (
            .in0(N__48154),
            .in1(N__45882),
            .in2(_gnd_net_),
            .in3(N__45927),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_21_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_21_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_21_11_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_21_11_1  (
            .in0(N__45862),
            .in1(N__45841),
            .in2(_gnd_net_),
            .in3(N__48149),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_21_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_21_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_21_11_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_21_11_6  (
            .in0(N__48150),
            .in1(N__45788),
            .in2(_gnd_net_),
            .in3(N__45769),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_21_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_21_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_21_12_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_24_LC_21_12_2  (
            .in0(N__45858),
            .in1(N__45830),
            .in2(_gnd_net_),
            .in3(N__48202),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47683),
            .ce(N__47236),
            .sr(N__46820));
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_21_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_21_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_21_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_26_LC_21_12_5  (
            .in0(N__48201),
            .in1(N__45786),
            .in2(_gnd_net_),
            .in3(N__45756),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47683),
            .ce(N__47236),
            .sr(N__46820));
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_21_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_21_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_21_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_27_LC_21_12_6  (
            .in0(N__48287),
            .in1(N__48227),
            .in2(_gnd_net_),
            .in3(N__48203),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47683),
            .ce(N__47236),
            .sr(N__46820));
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_21_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_21_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_21_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_25_LC_21_12_7  (
            .in0(N__48200),
            .in1(N__47762),
            .in2(_gnd_net_),
            .in3(N__47718),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47683),
            .ce(N__47236),
            .sr(N__46820));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_21_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_21_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_21_13_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_21_13_0  (
            .in0(N__46445),
            .in1(N__46435),
            .in2(N__46414),
            .in3(N__46388),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_21_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_21_13_4 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_21_13_4  (
            .in0(N__46444),
            .in1(N__46436),
            .in2(N__46415),
            .in3(N__46387),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_21_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_21_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_21_13_7 .LUT_INIT=16'b1101111100001101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_21_13_7  (
            .in0(N__46366),
            .in1(N__46345),
            .in2(N__46334),
            .in3(N__46306),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_1 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_1  (
            .in0(N__46270),
            .in1(N__46209),
            .in2(_gnd_net_),
            .in3(N__46079),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MAIN
